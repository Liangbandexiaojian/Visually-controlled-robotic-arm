
// Efinity Top-level template
// Version: 2023.2.307.5.10
// Date: 2024-11-11 18:32

// Copyright (C) 2013 - 2023 Efinix Inc. All rights reserved.

// This file may be used as a starting point for Efinity synthesis top-level target.
// The port list here matches what is expected by Efinity constraint files generated
// by the Efinity Interface Designer.

// To use this:
//     #1)  Save this file with a different name to a different directory, where source files are kept.
//              Example: you may wish to save as D:\code\learning\a241111_03\Efinity\T35_Sensor_DDR3_LCD_Test.v
//     #2)  Add the newly saved file into Efinity project as design file
//     #3)  Edit the top level entity in Efinity project to:  T35_Sensor_DDR3_LCD_Test
//     #4)  Insert design content.


module T35_Sensor_DDR3_LCD_Test
(
  input AxiPllClkIn,
  input DdrPllClkIn,
  input key0,
  input [1:0] PllLocked,
  input hdmi_lock_i,
  input mipi_lock_i,
  input mipi0_scl_i,
  input mipi0_sda_i,
  input mipi1_scl_i,
  input mipi1_sda_i,
  input cmos_ctl0_i,
  input cmos_ctl1_i,
  input cmos_ctl2_i,
  input cmos_ctl3_i,
  input [7:0] cmos_data,
  input cmos_href,
  input cmos_sdat_IN,
  input cmos_vsync,
  input [3:0] mipi_rx_0_CNT_i,
  input [63:0] mipi_rx_0_DATA_i,
  input [17:0] mipi_rx_0_ERROR,
  input [3:0] mipi_rx_0_HSYNC_i,
  input [5:0] mipi_rx_0_TYPE_i,
  input [3:0] mipi_rx_0_ULPS,
  input mipi_rx_0_ULPS_CLK,
  input mipi_rx_0_VALID_i,
  input [1:0] mipi_rx_0_VC_i,
  input [3:0] mipi_rx_0_VSYNC_i,
  input [3:0] mipi_rx_1_CNT_i,
  input [63:0] mipi_rx_1_DATA_i,
  input [17:0] mipi_rx_1_ERROR,
  input [3:0] mipi_rx_1_HSYNC_i,
  input [5:0] mipi_rx_1_TYPE_i,
  input [3:0] mipi_rx_1_ULPS,
  input mipi_rx_1_ULPS_CLK,
  input mipi_rx_1_VALID_i,
  input [1:0] mipi_rx_1_VC_i,
  input [3:0] mipi_rx_1_VSYNC_i,
  input cmos_pclk,
  input mipi_clkcal_i,
  input mipi_pixclk_i,
  input mipi_clkesc_i,
  input Axi0Clk,
  input tx_slowclk,
  input tx_fastclk,
  input hdmi_clk2x_i,
  input hdmi_clk5x_i,
  input clk_cmos,
  input hdmi_clk1x_i,
  input jtag_inst1_CAPTURE,
  input jtag_inst1_DRCK,
  input jtag_inst1_RESET,
  input jtag_inst1_RUNTEST,
  input jtag_inst1_SEL,
  input jtag_inst1_SHIFT,
  input jtag_inst1_TCK,
  input jtag_inst1_TDI,
  input jtag_inst1_TMS,
  input jtag_inst1_UPDATE,
  input DdrCtrl_AREADY_0,
  input [7:0] DdrCtrl_BID_0,
  input DdrCtrl_BVALID_0,
  input [127:0] DdrCtrl_RDATA_0,
  input [7:0] DdrCtrl_RID_0,
  input DdrCtrl_RLAST_0,
  input [1:0] DdrCtrl_RRESP_0,
  input DdrCtrl_RVALID_0,
  input DdrCtrl_WREADY_0,
  output [7:0] led_data,
  output hdmi_resetn_o,
  output mipi_resetn_o,
  output lcd_pwm,
  output mipi0_scl_o,
  output mipi0_scl_oe,
  output mipi0_sda_o,
  output mipi0_sda_oe,
  output mipi1_scl_o,
  output mipi1_scl_oe,
  output mipi1_sda_o,
  output mipi1_sda_oe,
  output [1:0] mipi_trig_o,
  output zone_bit0,
  output zone_bit1,
  output zone_bit2,
  output [4:0] hdmi_tx0_o,
  output [4:0] hdmi_tx1_o,
  output [4:0] hdmi_tx2_o,
  output [4:0] hdmi_txc_o,
  output [6:0] lvds_tx0_DATA,
  output [6:0] lvds_tx1_DATA,
  output [6:0] lvds_tx2_DATA,
  output [6:0] lvds_tx3_DATA,
  output [6:0] lvds_tx_clk_DATA,
  output cmos_ctl0_o,
  output cmos_ctl0_oe,
  output cmos_ctl1_o,
  output cmos_ctl1_oe,
  output cmos_ctl2_o,
  output cmos_ctl2_oe,
  output cmos_ctl3_o,
  output cmos_ctl3_oe,
  output cmos_sclk,
  output cmos_sdat_OUT,
  output cmos_sdat_OE,
  output mipi_rx_0_CLEAR,
  output mipi_rx_0_DPHY_RSTN_o,
  output [1:0] mipi_rx_0_LANES_o,
  output mipi_rx_0_RSTN_o,
  output [3:0] mipi_rx_0_VC_ENA_o,
  output mipi_rx_1_CLEAR,
  output mipi_rx_1_DPHY_RSTN_o,
  output [1:0] mipi_rx_1_LANES_o,
  output mipi_rx_1_RSTN_o,
  output [3:0] mipi_rx_1_VC_ENA_o,
  output jtag_inst1_TDO,
  output [31:0] DdrCtrl_AADDR_0,
  output [1:0] DdrCtrl_ABURST_0,
  output [7:0] DdrCtrl_AID_0,
  output [7:0] DdrCtrl_ALEN_0,
  output [1:0] DdrCtrl_ALOCK_0,
  output [2:0] DdrCtrl_ASIZE_0,
  output DdrCtrl_ATYPE_0,
  output DdrCtrl_AVALID_0,
  output DdrCtrl_BREADY_0,
  output DdrCtrl_CFG_SEQ_RST,
  output DdrCtrl_CFG_SEQ_START,
  output DdrCtrl_RREADY_0,
  output DdrCtrl_RSTN,
  output [127:0] DdrCtrl_WDATA_0,
  output [7:0] DdrCtrl_WID_0,
  output DdrCtrl_WLAST_0,
  output [15:0] DdrCtrl_WSTRB_0,
  output DdrCtrl_WVALID_0
);


endmodule

