
//
// Verific Verilog Description of module T35_Sensor_DDR3_LCD_Test
//

module T35_Sensor_DDR3_LCD_Test (AxiPllClkIn, DdrPllClkIn, Axi0Clk, hdmi_resetn_o, 
            mipi_resetn_o, mipi_clkcal_i, mipi_clkesc_i, mipi_pixclk_i, 
            hdmi_clk1x_i, hdmi_clk2x_i, hdmi_clk5x_i, clk_cmos, tx_slowclk, 
            tx_fastclk, PllLocked, hdmi_lock_i, mipi_lock_i, DdrCtrl_RSTN, 
            DdrCtrl_CFG_SEQ_RST, DdrCtrl_CFG_SEQ_START, DdrCtrl_AID_0, 
            DdrCtrl_AADDR_0, DdrCtrl_ALEN_0, DdrCtrl_ASIZE_0, DdrCtrl_ABURST_0, 
            DdrCtrl_ALOCK_0, DdrCtrl_AVALID_0, DdrCtrl_AREADY_0, DdrCtrl_ATYPE_0, 
            DdrCtrl_WID_0, DdrCtrl_WDATA_0, DdrCtrl_WSTRB_0, DdrCtrl_WLAST_0, 
            DdrCtrl_WVALID_0, DdrCtrl_WREADY_0, DdrCtrl_RID_0, DdrCtrl_RDATA_0, 
            DdrCtrl_RLAST_0, DdrCtrl_RVALID_0, DdrCtrl_RREADY_0, DdrCtrl_RRESP_0, 
            DdrCtrl_BID_0, DdrCtrl_BVALID_0, DdrCtrl_BREADY_0, led_data, 
            lcd_pwm, lvds_tx_clk_DATA, lvds_tx0_DATA, lvds_tx1_DATA, 
            lvds_tx2_DATA, lvds_tx3_DATA, hdmi_tx0_o, hdmi_tx1_o, hdmi_tx2_o, 
            hdmi_txc_o, zone_bit0, zone_bit1, zone_bit2, key0, cmos_pclk, 
            cmos_vsync, cmos_href, cmos_data, cmos_sclk, cmos_sdat_IN, 
            cmos_sdat_OUT, cmos_sdat_OE, mipi0_scl_i, mipi0_scl_o, mipi0_scl_oe, 
            mipi0_sda_i, mipi0_sda_o, mipi0_sda_oe, mipi1_scl_i, mipi1_scl_o, 
            mipi1_scl_oe, mipi1_sda_i, mipi1_sda_o, mipi1_sda_oe, mipi_trig_o, 
            mipi_rx_0_RSTN_o, mipi_rx_0_DPHY_RSTN_o, mipi_rx_0_VC_ENA_o, 
            mipi_rx_0_LANES_o, mipi_rx_1_RSTN_o, mipi_rx_1_DPHY_RSTN_o, 
            mipi_rx_1_VC_ENA_o, mipi_rx_1_LANES_o, mipi_rx_0_VC_i, mipi_rx_0_VSYNC_i, 
            mipi_rx_0_HSYNC_i, mipi_rx_0_DATA_i, mipi_rx_0_CNT_i, mipi_rx_0_TYPE_i, 
            mipi_rx_0_VALID_i, mipi_rx_1_VC_i, mipi_rx_1_VSYNC_i, mipi_rx_1_HSYNC_i, 
            mipi_rx_1_DATA_i, mipi_rx_1_CNT_i, mipi_rx_1_TYPE_i, mipi_rx_1_VALID_i, 
            mipi_rx_0_ULPS, mipi_rx_0_ULPS_CLK, mipi_rx_0_CLEAR, mipi_rx_0_ERROR, 
            mipi_rx_1_ULPS, mipi_rx_1_ULPS_CLK, mipi_rx_1_CLEAR, mipi_rx_1_ERROR);
    input AxiPllClkIn /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrPllClkIn /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input Axi0Clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output hdmi_resetn_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_resetn_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input mipi_clkcal_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_clkesc_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_pixclk_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk1x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk2x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk5x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input clk_cmos /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_slowclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_fastclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [1:0]PllLocked /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_lock_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_lock_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_RST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_START /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_AID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [31:0]DdrCtrl_AADDR_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_ALEN_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [2:0]DdrCtrl_ASIZE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ABURST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ALOCK_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_AVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_AREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_ATYPE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_WID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [127:0]DdrCtrl_WDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]DdrCtrl_WSTRB_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_WREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_RID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [127:0]DdrCtrl_RDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_RREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]DdrCtrl_RRESP_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_BID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_BVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_BREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]led_data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output lcd_pwm /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx_clk_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx0_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx1_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx2_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx3_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx0_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx1_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx2_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_txc_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output zone_bit0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output zone_bit1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output zone_bit2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input key0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input cmos_pclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input cmos_vsync /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input cmos_href /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]cmos_data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_sclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_sdat_IN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_sdat_OUT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output cmos_sdat_OE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input mipi0_scl_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi0_scl_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi0_scl_oe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input mipi0_sda_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi0_sda_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi0_sda_oe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input mipi1_scl_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi1_scl_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi1_scl_oe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input mipi1_sda_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi1_sda_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi1_sda_oe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]mipi_trig_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_rx_0_RSTN_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_rx_0_DPHY_RSTN_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]mipi_rx_0_VC_ENA_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]mipi_rx_0_LANES_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_rx_1_RSTN_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_rx_1_DPHY_RSTN_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]mipi_rx_1_VC_ENA_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]mipi_rx_1_LANES_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]mipi_rx_0_VC_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_0_VSYNC_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_0_HSYNC_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [63:0]mipi_rx_0_DATA_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_0_CNT_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [5:0]mipi_rx_0_TYPE_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_rx_0_VALID_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [1:0]mipi_rx_1_VC_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_1_VSYNC_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_1_HSYNC_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [63:0]mipi_rx_1_DATA_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_1_CNT_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [5:0]mipi_rx_1_TYPE_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_rx_1_VALID_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_0_ULPS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_rx_0_ULPS_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi_rx_0_CLEAR /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [17:0]mipi_rx_0_ERROR /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_rx_1_ULPS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_rx_1_ULPS_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi_rx_1_CLEAR /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [17:0]mipi_rx_1_ERROR /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire n927_2;
    wire n938_2;
    wire n949_2;
    wire n33_2;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire n926_2;
    wire n925_2;
    wire n924_2;
    wire n923_2;
    wire n937_2;
    wire n936_2;
    wire n935_2;
    wire n934_2;
    wire n948_2;
    wire n947_2;
    wire n946_2;
    wire n945_2;
    wire n32_2;
    wire n31_2;
    wire n30_2;
    wire n29_2;
    wire n28_2;
    wire n27_2;
    wire n26_2;
    
    wire \Axi0ResetReg[2] , n405, n406, \ResetShiftReg[0] , r_XYCrop0_frame_vsync, 
        \r_XYCrop0_frame_Gray[0] , r_XYCrop0_frame_href, r_XYCrop0_frame_de, 
        r_hdmi_rst_n, rc_hdmi_tx, n419, n420, n421, \PowerOnResetCnt[0] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] , 
        n431, n432, \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] , n453, n454, \u_i2c_timing_ctrl_16bit/clk_cnt[0] , 
        n456, n457, \u_i2c_timing_ctrl_16bit/current_state[0] , \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk , 
        \u_i2c_timing_ctrl_16bit/i2c_transfer_en , \i2c_config_index[0] , 
        n463, n464, \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] , \u_i2c_timing_ctrl_16bit/i2c_wdata[0] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[1] , \u_i2c_timing_ctrl_16bit/delay_cnt[0] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[1] , \u_i2c_timing_ctrl_16bit/clk_cnt[2] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[3] , \u_i2c_timing_ctrl_16bit/clk_cnt[4] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[5] , \u_i2c_timing_ctrl_16bit/clk_cnt[6] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[7] , \u_i2c_timing_ctrl_16bit/clk_cnt[8] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[9] , \u_i2c_timing_ctrl_16bit/clk_cnt[10] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[11] , \u_i2c_timing_ctrl_16bit/clk_cnt[12] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[13] , \u_i2c_timing_ctrl_16bit/clk_cnt[14] , 
        \u_i2c_timing_ctrl_16bit/clk_cnt[15] , \u_i2c_timing_ctrl_16bit/current_state[1] , 
        \u_i2c_timing_ctrl_16bit/current_state[2] , \u_i2c_timing_ctrl_16bit/current_state[3] , 
        \i2c_config_index[1] , \i2c_config_index[2] , \i2c_config_index[3] , 
        \i2c_config_index[4] , \i2c_config_index[5] , \i2c_config_index[6] , 
        \i2c_config_index[7] , \i2c_config_index[8] , n501, n502, \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] , 
        \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2] , \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3] , 
        \u_i2c_timing_ctrl_16bit/i2c_wdata[1] , \u_i2c_timing_ctrl_16bit/i2c_wdata[2] , 
        \u_i2c_timing_ctrl_16bit/i2c_wdata[3] , \u_i2c_timing_ctrl_16bit/i2c_wdata[4] , 
        \u_i2c_timing_ctrl_16bit/i2c_wdata[5] , \u_i2c_timing_ctrl_16bit/i2c_wdata[6] , 
        \u_i2c_timing_ctrl_16bit/i2c_wdata[7] , \u_i2c_timing_ctrl_16bit/delay_cnt[2] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[3] , \u_i2c_timing_ctrl_16bit/delay_cnt[4] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[5] , \u_i2c_timing_ctrl_16bit/delay_cnt[6] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[7] , \u_i2c_timing_ctrl_16bit/delay_cnt[8] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[9] , \u_i2c_timing_ctrl_16bit/delay_cnt[10] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[11] , \u_i2c_timing_ctrl_16bit/delay_cnt[12] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[13] , \u_i2c_timing_ctrl_16bit/delay_cnt[14] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[15] , \u_i2c_timing_ctrl_16bit/delay_cnt[16] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[17] , \u_i2c_timing_ctrl_16bit/delay_cnt[18] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[19] , \u_i2c_timing_ctrl_16bit/delay_cnt[20] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[21] , \u_i2c_timing_ctrl_16bit/delay_cnt[22] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[23] , \u_i2c_timing_ctrl_16bit/delay_cnt[24] , 
        \u_i2c_timing_ctrl_16bit/delay_cnt[25] , \u_i2c_timing_ctrl_16bit/delay_cnt[26] , 
        \u_Sensor_Image_XYCrop_0/image_ypos[11] , \u_Sensor_Image_XYCrop_0/image_ypos[10] , 
        \u_Sensor_Image_XYCrop_0/image_ypos[9] , n541, n542, \u_Sensor_Image_XYCrop_0/image_in_href_r , 
        \u_Sensor_Image_XYCrop_0/image_ypos[0] , n546, n547, \u_Sensor_Image_XYCrop_0/image_ypos[8] , 
        \u_Sensor_Image_XYCrop_0/image_ypos[7] , \w_XYCrop0_frame_Gray[5] , 
        \u_Sensor_Image_XYCrop_0/image_ypos[6] , \u_Sensor_Image_XYCrop_0/image_ypos[5] , 
        \u_Sensor_Image_XYCrop_0/image_xpos[0] , \w_XYCrop0_frame_Gray[3] , 
        \u_Sensor_Image_XYCrop_0/image_ypos[4] , \u_Sensor_Image_XYCrop_0/image_ypos[3] , 
        \w_XYCrop0_frame_Gray[4] , \u_Sensor_Image_XYCrop_0/image_ypos[2] , 
        \u_Sensor_Image_XYCrop_0/image_ypos[1] , \w_XYCrop0_frame_Gray[6] , 
        \w_XYCrop0_frame_Gray[7] , \w_XYCrop0_frame_Gray[2] , \w_XYCrop0_frame_Gray[1] , 
        \u_Sensor_Image_XYCrop_0/image_xpos[1] , \u_Sensor_Image_XYCrop_0/image_xpos[2] , 
        \u_Sensor_Image_XYCrop_0/image_xpos[3] , \u_Sensor_Image_XYCrop_0/image_xpos[4] , 
        \u_Sensor_Image_XYCrop_0/image_xpos[5] , \u_Sensor_Image_XYCrop_0/image_xpos[6] , 
        \u_Sensor_Image_XYCrop_0/image_xpos[7] , \u_Sensor_Image_XYCrop_0/image_xpos[8] , 
        \u_Sensor_Image_XYCrop_0/image_xpos[9] , \u_Sensor_Image_XYCrop_0/image_xpos[10] , 
        \u_Sensor_Image_XYCrop_0/image_xpos[11] , \r_XYCrop0_frame_Gray[1] , 
        \r_XYCrop0_frame_Gray[2] , \r_XYCrop0_frame_Gray[3] , \r_XYCrop0_frame_Gray[4] , 
        \r_XYCrop0_frame_Gray[5] , \r_XYCrop0_frame_Gray[6] , \r_XYCrop0_frame_Gray[7] , 
        \axi4_awar_mux/rs_req[0] , DdrCtrl_AWREADY_0, DdrCtrl_ARREADY_0, 
        \axi4_awar_mux/rs_req[1] , \u_axi4_ctrl_0/r_wframe_index_last[1] , 
        \DdrCtrl_ARADDR_0[23] , \DdrCtrl_ARADDR_0[22] , \u_axi4_ctrl_0/r_wframe_index_last[0] , 
        \u_axi4_ctrl_0/rs_w[0] , \DdrCtrl_AWADDR_0[0] , \u_axi4_ctrl_0/r_wframe_sync[0] , 
        \u_axi4_ctrl_0/rc_w_eof[0] , DdrCtrl_AWVALID_0, \u_axi4_ctrl_0/rc_burst[0] , 
        \u_axi4_ctrl_0/r_weof_pending , \u_axi4_ctrl_0/r_wframe_inc , \u_axi4_ctrl_0/rc_wfifo_we[0] , 
        \u_axi4_ctrl_0/rframe_vsync_dly , \u_axi4_ctrl_0/rfifo_cnt[1] , 
        \u_axi4_ctrl_0/rfifo_cnt[0] , \u_axi4_ctrl_0/rfifo_rst , n631, 
        n632, \u_axi4_ctrl_0/r_rfifo_rst , \u_axi4_ctrl_0/rc_rfifo_rd[0] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0] , \u_axi4_ctrl_0/r_rframe_inc , 
        \u_axi4_ctrl_0/rd_state.S_READ_IDLE , \u_axi4_ctrl_0/rd_state.S_READ_ADDR , 
        \u_axi4_ctrl_0/rd_state.S_READ_DATA , DdrCtrl_ARVALID_0, \u_axi4_ctrl_0/r_rd_pend , 
        \u_axi4_ctrl_0/rfifo_wenb , \u_axi4_ctrl_0/rfifo_wdata[3] , \u_axi4_ctrl_0/rfifo_wdata[2] , 
        \u_axi4_ctrl_0/rfifo_wdata[1] , \u_axi4_ctrl_0/rfifo_wdata[0] , 
        \u_axi4_ctrl_0/rs_w[1] , \DdrCtrl_AWADDR_0[22] , \DdrCtrl_AWADDR_0[1] , 
        \DdrCtrl_AWADDR_0[2] , \DdrCtrl_AWADDR_0[3] , \DdrCtrl_AWADDR_0[4] , 
        \DdrCtrl_AWADDR_0[5] , \DdrCtrl_AWADDR_0[6] , \DdrCtrl_AWADDR_0[7] , 
        \DdrCtrl_AWADDR_0[8] , \DdrCtrl_AWADDR_0[9] , \DdrCtrl_AWADDR_0[10] , 
        \DdrCtrl_AWADDR_0[11] , \DdrCtrl_AWADDR_0[12] , \DdrCtrl_AWADDR_0[13] , 
        \DdrCtrl_AWADDR_0[14] , \DdrCtrl_AWADDR_0[15] , \DdrCtrl_AWADDR_0[16] , 
        \DdrCtrl_AWADDR_0[17] , \DdrCtrl_AWADDR_0[18] , \DdrCtrl_AWADDR_0[19] , 
        \DdrCtrl_AWADDR_0[20] , \DdrCtrl_AWADDR_0[21] , \u_axi4_ctrl_0/r_wframe_sync[1] , 
        \u_axi4_ctrl_0/rc_burst[1] , \u_axi4_ctrl_0/rc_burst[2] , \u_axi4_ctrl_0/rc_burst[3] , 
        \u_axi4_ctrl_0/rc_burst[4] , \u_axi4_ctrl_0/rc_burst[5] , \u_axi4_ctrl_0/rc_burst[6] , 
        \u_axi4_ctrl_0/rc_burst[7] , \u_axi4_ctrl_0/r_wfifo_wdata[8] , \u_axi4_ctrl_0/r_wfifo_wdata[9] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[10] , \u_axi4_ctrl_0/r_wfifo_wdata[11] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[12] , \u_axi4_ctrl_0/r_wfifo_wdata[13] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[14] , \u_axi4_ctrl_0/r_wfifo_wdata[15] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[16] , \u_axi4_ctrl_0/r_wfifo_wdata[17] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[18] , \u_axi4_ctrl_0/r_wfifo_wdata[19] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[20] , \u_axi4_ctrl_0/r_wfifo_wdata[21] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[22] , \u_axi4_ctrl_0/r_wfifo_wdata[23] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[24] , \u_axi4_ctrl_0/r_wfifo_wdata[25] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[26] , \u_axi4_ctrl_0/r_wfifo_wdata[27] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[28] , \u_axi4_ctrl_0/r_wfifo_wdata[29] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[30] , \u_axi4_ctrl_0/r_wfifo_wdata[31] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[32] , \u_axi4_ctrl_0/r_wfifo_wdata[33] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[34] , \u_axi4_ctrl_0/r_wfifo_wdata[35] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[36] , \u_axi4_ctrl_0/r_wfifo_wdata[37] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[38] , \u_axi4_ctrl_0/r_wfifo_wdata[39] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[40] , \u_axi4_ctrl_0/r_wfifo_wdata[41] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[42] , \u_axi4_ctrl_0/r_wfifo_wdata[43] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[44] , \u_axi4_ctrl_0/r_wfifo_wdata[45] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[46] , \u_axi4_ctrl_0/r_wfifo_wdata[47] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[48] , \u_axi4_ctrl_0/r_wfifo_wdata[49] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[50] , \u_axi4_ctrl_0/r_wfifo_wdata[51] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[52] , \u_axi4_ctrl_0/r_wfifo_wdata[53] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[54] , \u_axi4_ctrl_0/r_wfifo_wdata[55] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[56] , \u_axi4_ctrl_0/r_wfifo_wdata[57] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[58] , \u_axi4_ctrl_0/r_wfifo_wdata[59] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[60] , \u_axi4_ctrl_0/r_wfifo_wdata[61] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[62] , \u_axi4_ctrl_0/r_wfifo_wdata[63] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[64] , \u_axi4_ctrl_0/r_wfifo_wdata[65] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[66] , \u_axi4_ctrl_0/r_wfifo_wdata[67] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[68] , \u_axi4_ctrl_0/r_wfifo_wdata[69] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[70] , \u_axi4_ctrl_0/r_wfifo_wdata[71] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[72] , \u_axi4_ctrl_0/r_wfifo_wdata[73] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[74] , \u_axi4_ctrl_0/r_wfifo_wdata[75] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[76] , \u_axi4_ctrl_0/r_wfifo_wdata[77] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[78] , \u_axi4_ctrl_0/r_wfifo_wdata[79] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[80] , \u_axi4_ctrl_0/r_wfifo_wdata[81] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[82] , \u_axi4_ctrl_0/r_wfifo_wdata[83] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[84] , \u_axi4_ctrl_0/r_wfifo_wdata[85] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[86] , \u_axi4_ctrl_0/r_wfifo_wdata[87] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[88] , \u_axi4_ctrl_0/r_wfifo_wdata[89] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[90] , \u_axi4_ctrl_0/r_wfifo_wdata[91] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[92] , \u_axi4_ctrl_0/r_wfifo_wdata[93] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[94] , \u_axi4_ctrl_0/r_wfifo_wdata[95] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[96] , \u_axi4_ctrl_0/r_wfifo_wdata[97] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[98] , \u_axi4_ctrl_0/r_wfifo_wdata[99] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[100] , \u_axi4_ctrl_0/r_wfifo_wdata[101] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[102] , \u_axi4_ctrl_0/r_wfifo_wdata[103] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[104] , \u_axi4_ctrl_0/r_wfifo_wdata[105] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[106] , \u_axi4_ctrl_0/r_wfifo_wdata[107] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[108] , \u_axi4_ctrl_0/r_wfifo_wdata[109] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[110] , \u_axi4_ctrl_0/r_wfifo_wdata[111] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[112] , \u_axi4_ctrl_0/r_wfifo_wdata[113] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[114] , \u_axi4_ctrl_0/r_wfifo_wdata[115] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[116] , \u_axi4_ctrl_0/r_wfifo_wdata[117] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[118] , \u_axi4_ctrl_0/r_wfifo_wdata[119] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[120] , \u_axi4_ctrl_0/r_wfifo_wdata[121] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[122] , \u_axi4_ctrl_0/r_wfifo_wdata[123] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[124] , \u_axi4_ctrl_0/r_wfifo_wdata[125] , 
        \u_axi4_ctrl_0/r_wfifo_wdata[126] , \u_axi4_ctrl_0/r_wfifo_wdata[127] , 
        \u_axi4_ctrl_0/rc_wfifo_we[1] , \u_axi4_ctrl_0/rc_wfifo_we[2] , 
        \u_axi4_ctrl_0/rc_wfifo_we[3] , n929, n930, \u_axi4_ctrl_0/w_rframe_data_gen[48] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[49] , \u_axi4_ctrl_0/w_rframe_data_gen[50] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[51] , \u_axi4_ctrl_0/w_rframe_data_gen[52] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[53] , \u_axi4_ctrl_0/w_rframe_data_gen[54] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[55] , \u_axi4_ctrl_0/w_rframe_data_gen[56] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[57] , \u_axi4_ctrl_0/w_rframe_data_gen[58] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[59] , \u_axi4_ctrl_0/w_rframe_data_gen[60] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[61] , \u_axi4_ctrl_0/w_rframe_data_gen[62] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[63] , \u_axi4_ctrl_0/w_rframe_data_gen[64] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[65] , \u_axi4_ctrl_0/w_rframe_data_gen[66] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[67] , n954, n955, \u_axi4_ctrl_0/w_wfifo_empty , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] , n958, n959, 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] , n961, n962, 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] , 
        n977, n978, n979, \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        \u_axi4_ctrl_0/rfifo_cnt[2] , \u_axi4_ctrl_0/rfifo_cnt[3] , \u_axi4_ctrl_0/rfifo_cnt[4] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[0] , \u_axi4_ctrl_0/w_rframe_data_gen[1] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[2] , \u_axi4_ctrl_0/w_rframe_data_gen[3] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[4] , \u_axi4_ctrl_0/w_rframe_data_gen[5] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[6] , \u_axi4_ctrl_0/w_rframe_data_gen[7] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[8] , \u_axi4_ctrl_0/w_rframe_data_gen[9] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[10] , \u_axi4_ctrl_0/w_rframe_data_gen[11] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[12] , \u_axi4_ctrl_0/w_rframe_data_gen[13] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[14] , \u_axi4_ctrl_0/w_rframe_data_gen[15] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[108] , \u_axi4_ctrl_0/w_rframe_data_gen[109] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[110] , \u_axi4_ctrl_0/w_rframe_data_gen[111] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[112] , \u_axi4_ctrl_0/w_rframe_data_gen[113] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[114] , \u_axi4_ctrl_0/w_rframe_data_gen[115] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[116] , \u_axi4_ctrl_0/w_rframe_data_gen[117] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[118] , \u_axi4_ctrl_0/w_rframe_data_gen[119] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[120] , \u_axi4_ctrl_0/w_rframe_data_gen[121] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[122] , \u_axi4_ctrl_0/w_rframe_data_gen[123] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[124] , \u_axi4_ctrl_0/w_rframe_data_gen[125] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[126] , \u_axi4_ctrl_0/w_rframe_data_gen[127] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[16] , \u_axi4_ctrl_0/w_rframe_data_gen[17] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[18] , \u_axi4_ctrl_0/w_rframe_data_gen[19] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[20] , \u_axi4_ctrl_0/w_rframe_data_gen[21] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[22] , \u_axi4_ctrl_0/w_rframe_data_gen[23] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[24] , \u_axi4_ctrl_0/w_rframe_data_gen[25] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[26] , \u_axi4_ctrl_0/w_rframe_data_gen[27] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[28] , \u_axi4_ctrl_0/w_rframe_data_gen[29] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[30] , \u_axi4_ctrl_0/w_rframe_data_gen[31] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[68] , \u_axi4_ctrl_0/w_rframe_data_gen[69] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[70] , \u_axi4_ctrl_0/w_rframe_data_gen[71] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[72] , \u_axi4_ctrl_0/w_rframe_data_gen[73] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[74] , \u_axi4_ctrl_0/w_rframe_data_gen[75] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[76] , \u_axi4_ctrl_0/w_rframe_data_gen[77] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[78] , \u_axi4_ctrl_0/w_rframe_data_gen[79] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[80] , \u_axi4_ctrl_0/w_rframe_data_gen[81] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[82] , \u_axi4_ctrl_0/w_rframe_data_gen[83] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[84] , \u_axi4_ctrl_0/w_rframe_data_gen[85] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[86] , \u_axi4_ctrl_0/w_rframe_data_gen[87] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[88] , \u_axi4_ctrl_0/w_rframe_data_gen[89] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[90] , \u_axi4_ctrl_0/w_rframe_data_gen[91] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[92] , \u_axi4_ctrl_0/w_rframe_data_gen[93] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[94] , \u_axi4_ctrl_0/w_rframe_data_gen[95] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[96] , \u_axi4_ctrl_0/w_rframe_data_gen[97] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[98] , \u_axi4_ctrl_0/w_rframe_data_gen[99] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[100] , \u_axi4_ctrl_0/w_rframe_data_gen[101] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[102] , \u_axi4_ctrl_0/w_rframe_data_gen[103] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[104] , \u_axi4_ctrl_0/w_rframe_data_gen[105] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[106] , \u_axi4_ctrl_0/w_rframe_data_gen[107] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[32] , \u_axi4_ctrl_0/w_rframe_data_gen[33] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[34] , \u_axi4_ctrl_0/w_rframe_data_gen[35] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[36] , \u_axi4_ctrl_0/w_rframe_data_gen[37] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[38] , \u_axi4_ctrl_0/w_rframe_data_gen[39] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[40] , \u_axi4_ctrl_0/w_rframe_data_gen[41] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[42] , \u_axi4_ctrl_0/w_rframe_data_gen[43] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[44] , \u_axi4_ctrl_0/w_rframe_data_gen[45] , 
        \u_axi4_ctrl_0/w_rframe_data_gen[46] , \u_axi4_ctrl_0/w_rframe_data_gen[47] , 
        n1194, n1195, n1196, n1197, n1201, n1202, \u_axi4_ctrl_0/w_rfifo_empty , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] , n1205, n1206, 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] , n1208, n1209, 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] , 
        n1225, \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        \u_axi4_ctrl_0/rc_rfifo_rd[1] , \u_axi4_ctrl_0/rc_rfifo_rd[2] , 
        \lcd_data[0] , \lcd_data[1] , \lcd_data[2] , \lcd_data[3] , 
        \lcd_data[4] , \lcd_data[5] , \lcd_data[6] , \lcd_data[7] , 
        \lcd_data[8] , \lcd_data[9] , \lcd_data[10] , \lcd_data[11] , 
        \lcd_data[12] , \lcd_data[13] , \lcd_data[14] , \lcd_data[15] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[16] , \u_axi4_ctrl_0/r_rframe_data_gen[17] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[18] , \u_axi4_ctrl_0/r_rframe_data_gen[19] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[20] , \u_axi4_ctrl_0/r_rframe_data_gen[21] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[22] , \u_axi4_ctrl_0/r_rframe_data_gen[23] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[24] , \u_axi4_ctrl_0/r_rframe_data_gen[25] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[26] , \u_axi4_ctrl_0/r_rframe_data_gen[27] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[28] , \u_axi4_ctrl_0/r_rframe_data_gen[29] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[30] , \u_axi4_ctrl_0/r_rframe_data_gen[31] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[32] , \u_axi4_ctrl_0/r_rframe_data_gen[33] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[34] , \u_axi4_ctrl_0/r_rframe_data_gen[35] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[36] , \u_axi4_ctrl_0/r_rframe_data_gen[37] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[38] , \u_axi4_ctrl_0/r_rframe_data_gen[39] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[40] , \u_axi4_ctrl_0/r_rframe_data_gen[41] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[42] , \u_axi4_ctrl_0/r_rframe_data_gen[43] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[44] , \u_axi4_ctrl_0/r_rframe_data_gen[45] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[46] , \u_axi4_ctrl_0/r_rframe_data_gen[47] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[48] , \u_axi4_ctrl_0/r_rframe_data_gen[49] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[50] , \u_axi4_ctrl_0/r_rframe_data_gen[51] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[52] , \u_axi4_ctrl_0/r_rframe_data_gen[53] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[54] , \u_axi4_ctrl_0/r_rframe_data_gen[55] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[56] , \u_axi4_ctrl_0/r_rframe_data_gen[57] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[58] , \u_axi4_ctrl_0/r_rframe_data_gen[59] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[60] , \u_axi4_ctrl_0/r_rframe_data_gen[61] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[62] , \u_axi4_ctrl_0/r_rframe_data_gen[63] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[64] , \u_axi4_ctrl_0/r_rframe_data_gen[65] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[66] , \u_axi4_ctrl_0/r_rframe_data_gen[67] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[68] , \u_axi4_ctrl_0/r_rframe_data_gen[69] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[70] , \u_axi4_ctrl_0/r_rframe_data_gen[71] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[72] , \u_axi4_ctrl_0/r_rframe_data_gen[73] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[74] , \u_axi4_ctrl_0/r_rframe_data_gen[75] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[76] , \u_axi4_ctrl_0/r_rframe_data_gen[77] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[78] , \u_axi4_ctrl_0/r_rframe_data_gen[79] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[80] , \u_axi4_ctrl_0/r_rframe_data_gen[81] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[82] , \u_axi4_ctrl_0/r_rframe_data_gen[83] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[84] , \u_axi4_ctrl_0/r_rframe_data_gen[85] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[86] , \u_axi4_ctrl_0/r_rframe_data_gen[87] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[88] , \u_axi4_ctrl_0/r_rframe_data_gen[89] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[90] , \u_axi4_ctrl_0/r_rframe_data_gen[91] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[92] , \u_axi4_ctrl_0/r_rframe_data_gen[93] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[94] , \u_axi4_ctrl_0/r_rframe_data_gen[95] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[96] , \u_axi4_ctrl_0/r_rframe_data_gen[97] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[98] , \u_axi4_ctrl_0/r_rframe_data_gen[99] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[100] , \u_axi4_ctrl_0/r_rframe_data_gen[101] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[102] , \u_axi4_ctrl_0/r_rframe_data_gen[103] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[104] , \u_axi4_ctrl_0/r_rframe_data_gen[105] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[106] , \u_axi4_ctrl_0/r_rframe_data_gen[107] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[108] , \u_axi4_ctrl_0/r_rframe_data_gen[109] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[110] , \u_axi4_ctrl_0/r_rframe_data_gen[111] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[112] , \u_axi4_ctrl_0/r_rframe_data_gen[113] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[114] , \u_axi4_ctrl_0/r_rframe_data_gen[115] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[116] , \u_axi4_ctrl_0/r_rframe_data_gen[117] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[118] , \u_axi4_ctrl_0/r_rframe_data_gen[119] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[120] , \u_axi4_ctrl_0/r_rframe_data_gen[121] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[122] , \u_axi4_ctrl_0/r_rframe_data_gen[123] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[124] , \u_axi4_ctrl_0/r_rframe_data_gen[125] , 
        \u_axi4_ctrl_0/r_rframe_data_gen[126] , \u_axi4_ctrl_0/r_rframe_data_gen[127] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1] , \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3] , \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5] , \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7] , \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9] , \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11] , \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13] , \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14] , 
        \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15] , n1479, n1480, n617, 
        n618, n619, n620, n621, n622, n623, n624, n625, n626, 
        n627, n628, n629, \DdrCtrl_ARADDR_0[8] , \DdrCtrl_ARADDR_0[9] , 
        \DdrCtrl_ARADDR_0[10] , \DdrCtrl_ARADDR_0[11] , \DdrCtrl_ARADDR_0[12] , 
        \DdrCtrl_ARADDR_0[13] , \DdrCtrl_ARADDR_0[14] , \DdrCtrl_ARADDR_0[15] , 
        \DdrCtrl_ARADDR_0[16] , \DdrCtrl_ARADDR_0[17] , \DdrCtrl_ARADDR_0[18] , 
        \DdrCtrl_ARADDR_0[19] , \DdrCtrl_ARADDR_0[20] , \DdrCtrl_ARADDR_0[21] , 
        n682, n683, n684, n685, n686, n687, n688, n689, n690, 
        n691, n692, n693, n694, \u_axi4_ctrl_0/rfifo_wdata[4] , \u_axi4_ctrl_0/rfifo_wdata[5] , 
        \u_axi4_ctrl_0/rfifo_wdata[6] , \u_axi4_ctrl_0/rfifo_wdata[7] , 
        \u_axi4_ctrl_0/rfifo_wdata[8] , \u_axi4_ctrl_0/rfifo_wdata[9] , 
        \u_axi4_ctrl_0/rfifo_wdata[10] , \u_axi4_ctrl_0/rfifo_wdata[11] , 
        \u_axi4_ctrl_0/rfifo_wdata[12] , \u_axi4_ctrl_0/rfifo_wdata[13] , 
        \u_axi4_ctrl_0/rfifo_wdata[14] , \u_axi4_ctrl_0/rfifo_wdata[15] , 
        \u_axi4_ctrl_0/rfifo_wdata[16] , \u_axi4_ctrl_0/rfifo_wdata[17] , 
        \u_axi4_ctrl_0/rfifo_wdata[18] , \u_axi4_ctrl_0/rfifo_wdata[19] , 
        \u_axi4_ctrl_0/rfifo_wdata[20] , \u_axi4_ctrl_0/rfifo_wdata[21] , 
        \u_axi4_ctrl_0/rfifo_wdata[22] , \u_axi4_ctrl_0/rfifo_wdata[23] , 
        \u_axi4_ctrl_0/rfifo_wdata[24] , \u_axi4_ctrl_0/rfifo_wdata[25] , 
        \u_axi4_ctrl_0/rfifo_wdata[26] , \u_axi4_ctrl_0/rfifo_wdata[27] , 
        \u_axi4_ctrl_0/rfifo_wdata[28] , \u_axi4_ctrl_0/rfifo_wdata[29] , 
        \u_axi4_ctrl_0/rfifo_wdata[30] , \u_axi4_ctrl_0/rfifo_wdata[31] , 
        \u_axi4_ctrl_0/rfifo_wdata[32] , \u_axi4_ctrl_0/rfifo_wdata[33] , 
        \u_axi4_ctrl_0/rfifo_wdata[34] , \u_axi4_ctrl_0/rfifo_wdata[35] , 
        \u_axi4_ctrl_0/rfifo_wdata[36] , \u_axi4_ctrl_0/rfifo_wdata[37] , 
        \u_axi4_ctrl_0/rfifo_wdata[38] , \u_axi4_ctrl_0/rfifo_wdata[39] , 
        \u_axi4_ctrl_0/rfifo_wdata[40] , \u_axi4_ctrl_0/rfifo_wdata[41] , 
        \u_axi4_ctrl_0/rfifo_wdata[42] , \u_axi4_ctrl_0/rfifo_wdata[43] , 
        \u_axi4_ctrl_0/rfifo_wdata[44] , \u_axi4_ctrl_0/rfifo_wdata[45] , 
        \u_axi4_ctrl_0/rfifo_wdata[46] , \u_axi4_ctrl_0/rfifo_wdata[47] , 
        \u_axi4_ctrl_0/rfifo_wdata[48] , \u_axi4_ctrl_0/rfifo_wdata[49] , 
        \u_axi4_ctrl_0/rfifo_wdata[50] , \u_axi4_ctrl_0/rfifo_wdata[51] , 
        \u_axi4_ctrl_0/rfifo_wdata[52] , \u_axi4_ctrl_0/rfifo_wdata[53] , 
        \u_axi4_ctrl_0/rfifo_wdata[54] , \u_axi4_ctrl_0/rfifo_wdata[55] , 
        \u_axi4_ctrl_0/rfifo_wdata[56] , \u_axi4_ctrl_0/rfifo_wdata[57] , 
        \u_axi4_ctrl_0/rfifo_wdata[58] , \u_axi4_ctrl_0/rfifo_wdata[59] , 
        \u_axi4_ctrl_0/rfifo_wdata[60] , \u_axi4_ctrl_0/rfifo_wdata[61] , 
        \u_axi4_ctrl_0/rfifo_wdata[62] , \u_axi4_ctrl_0/rfifo_wdata[63] , 
        \u_axi4_ctrl_0/rfifo_wdata[64] , \u_axi4_ctrl_0/rfifo_wdata[65] , 
        \u_axi4_ctrl_0/rfifo_wdata[66] , \u_axi4_ctrl_0/rfifo_wdata[67] , 
        \u_axi4_ctrl_0/rfifo_wdata[68] , \u_axi4_ctrl_0/rfifo_wdata[69] , 
        \u_axi4_ctrl_0/rfifo_wdata[70] , \u_axi4_ctrl_0/rfifo_wdata[71] , 
        \u_axi4_ctrl_0/rfifo_wdata[72] , \u_axi4_ctrl_0/rfifo_wdata[73] , 
        \u_axi4_ctrl_0/rfifo_wdata[74] , \u_axi4_ctrl_0/rfifo_wdata[75] , 
        \u_axi4_ctrl_0/rfifo_wdata[76] , \u_axi4_ctrl_0/rfifo_wdata[77] , 
        \u_axi4_ctrl_0/rfifo_wdata[78] , \u_axi4_ctrl_0/rfifo_wdata[79] , 
        \u_axi4_ctrl_0/rfifo_wdata[80] , \u_axi4_ctrl_0/rfifo_wdata[81] , 
        \u_axi4_ctrl_0/rfifo_wdata[82] , \u_axi4_ctrl_0/rfifo_wdata[83] , 
        \u_axi4_ctrl_0/rfifo_wdata[84] , \u_axi4_ctrl_0/rfifo_wdata[85] , 
        \u_axi4_ctrl_0/rfifo_wdata[86] , \u_axi4_ctrl_0/rfifo_wdata[87] , 
        \u_axi4_ctrl_0/rfifo_wdata[88] , \u_axi4_ctrl_0/rfifo_wdata[89] , 
        \u_axi4_ctrl_0/rfifo_wdata[90] , \u_axi4_ctrl_0/rfifo_wdata[91] , 
        \u_axi4_ctrl_0/rfifo_wdata[92] , \u_axi4_ctrl_0/rfifo_wdata[93] , 
        \u_axi4_ctrl_0/rfifo_wdata[94] , \u_axi4_ctrl_0/rfifo_wdata[95] , 
        \u_axi4_ctrl_0/rfifo_wdata[96] , \u_axi4_ctrl_0/rfifo_wdata[97] , 
        \u_axi4_ctrl_0/rfifo_wdata[98] , \u_axi4_ctrl_0/rfifo_wdata[99] , 
        \u_axi4_ctrl_0/rfifo_wdata[100] , \u_axi4_ctrl_0/rfifo_wdata[101] , 
        \u_axi4_ctrl_0/rfifo_wdata[102] , \u_axi4_ctrl_0/rfifo_wdata[103] , 
        \u_axi4_ctrl_0/rfifo_wdata[104] , \u_axi4_ctrl_0/rfifo_wdata[105] , 
        \u_axi4_ctrl_0/rfifo_wdata[106] , \u_axi4_ctrl_0/rfifo_wdata[107] , 
        \u_axi4_ctrl_0/rfifo_wdata[108] , \u_axi4_ctrl_0/rfifo_wdata[109] , 
        \u_axi4_ctrl_0/rfifo_wdata[110] , \u_axi4_ctrl_0/rfifo_wdata[111] , 
        \u_axi4_ctrl_0/rfifo_wdata[112] , \u_axi4_ctrl_0/rfifo_wdata[113] , 
        \u_axi4_ctrl_0/rfifo_wdata[114] , \u_axi4_ctrl_0/rfifo_wdata[115] , 
        \u_axi4_ctrl_0/rfifo_wdata[116] , \u_axi4_ctrl_0/rfifo_wdata[117] , 
        \u_axi4_ctrl_0/rfifo_wdata[118] , \u_axi4_ctrl_0/rfifo_wdata[119] , 
        \u_axi4_ctrl_0/rfifo_wdata[120] , \u_axi4_ctrl_0/rfifo_wdata[121] , 
        \u_axi4_ctrl_0/rfifo_wdata[122] , \u_axi4_ctrl_0/rfifo_wdata[123] , 
        \u_axi4_ctrl_0/rfifo_wdata[124] , \u_axi4_ctrl_0/rfifo_wdata[125] , 
        \u_axi4_ctrl_0/rfifo_wdata[126] , \u_axi4_ctrl_0/rfifo_wdata[127] , 
        \DdrCtrl_AWADDR_0[23] , n1649, n1650, n1651, n1652, n1653, 
        n1654, \u_lcd_driver/vcnt[0] , lcd_hs, n1657, n1658, \u_lcd_driver/r_lcd_dv , 
        lcd_request, n1662, n1663, \lcd_xpos[0] , \lcd_ypos[0] , \u_lcd_driver/vcnt[1] , 
        \u_lcd_driver/vcnt[2] , \u_lcd_driver/vcnt[3] , \u_lcd_driver/vcnt[4] , 
        \u_lcd_driver/vcnt[5] , \u_lcd_driver/vcnt[6] , \u_lcd_driver/vcnt[7] , 
        \u_lcd_driver/vcnt[8] , \u_lcd_driver/vcnt[9] , \u_lcd_driver/vcnt[10] , 
        \u_lcd_driver/vcnt[11] , \u_lcd_driver/r_lcd_rgb[23] , n1679, 
        n1680, \lcd_xpos[1] , \lcd_xpos[2] , \lcd_xpos[3] , \lcd_xpos[4] , 
        \lcd_xpos[5] , \lcd_xpos[6] , \lcd_xpos[7] , \lcd_xpos[8] , 
        \lcd_xpos[9] , \lcd_xpos[10] , \lcd_xpos[11] , \lcd_ypos[1] , 
        \lcd_ypos[2] , \lcd_ypos[3] , \lcd_ypos[4] , \lcd_ypos[5] , 
        \lcd_ypos[6] , \lcd_ypos[7] , \lcd_ypos[8] , \lcd_ypos[9] , 
        \lcd_ypos[10] , \lcd_ypos[11] , \u_lcd_driver/hcnt[1] , \u_lcd_driver/hcnt[2] , 
        \u_lcd_driver/hcnt[3] , \u_lcd_driver/hcnt[4] , \u_lcd_driver/hcnt[5] , 
        \u_lcd_driver/hcnt[6] , \u_lcd_driver/hcnt[7] , \u_lcd_driver/hcnt[8] , 
        \u_lcd_driver/hcnt[9] , \u_lcd_driver/hcnt[10] , \u_lcd_driver/hcnt[11] , 
        n1714, n1715, n1716, n1717, \u_black_pixel_avg/y_sum[0] , 
        \u_black_pixel_avg/black_pixel_count[0] , n12161, \u_black_pixel_avg/x_sum[1] , 
        \u_black_pixel_avg/x_sum[0] , n1724, n1725, n1726, n1727, 
        n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
        n1736, n1737, n1738, \u_black_pixel_avg/y_sum[1] , \u_black_pixel_avg/y_sum[2] , 
        \u_black_pixel_avg/y_sum[3] , \u_black_pixel_avg/y_sum[4] , \u_black_pixel_avg/y_sum[5] , 
        \u_black_pixel_avg/y_sum[6] , \u_black_pixel_avg/y_sum[7] , \u_black_pixel_avg/y_sum[8] , 
        \u_black_pixel_avg/y_sum[9] , \u_black_pixel_avg/y_sum[10] , \u_black_pixel_avg/y_sum[11] , 
        \u_black_pixel_avg/y_sum[12] , \u_black_pixel_avg/y_sum[13] , \u_black_pixel_avg/y_sum[14] , 
        \u_black_pixel_avg/y_sum[15] , \u_black_pixel_avg/y_sum[16] , \u_black_pixel_avg/y_sum[17] , 
        \u_black_pixel_avg/y_sum[18] , \u_black_pixel_avg/y_sum[19] , \u_black_pixel_avg/y_sum[20] , 
        \u_black_pixel_avg/y_sum[21] , \u_black_pixel_avg/y_sum[22] , \u_black_pixel_avg/y_sum[23] , 
        \u_black_pixel_avg/y_sum[24] , \u_black_pixel_avg/y_sum[25] , \u_black_pixel_avg/y_sum[26] , 
        \u_black_pixel_avg/y_sum[27] , \u_black_pixel_avg/y_sum[28] , \u_black_pixel_avg/y_sum[29] , 
        \u_black_pixel_avg/y_sum[30] , \u_black_pixel_avg/y_sum[31] , \u_black_pixel_avg/black_pixel_count[1] , 
        \u_black_pixel_avg/black_pixel_count[2] , \u_black_pixel_avg/black_pixel_count[3] , 
        \u_black_pixel_avg/black_pixel_count[4] , \u_black_pixel_avg/black_pixel_count[5] , 
        \u_black_pixel_avg/black_pixel_count[6] , \u_black_pixel_avg/black_pixel_count[7] , 
        \u_black_pixel_avg/black_pixel_count[8] , \u_black_pixel_avg/black_pixel_count[9] , 
        \u_black_pixel_avg/black_pixel_count[10] , \u_black_pixel_avg/black_pixel_count[11] , 
        \u_black_pixel_avg/black_pixel_count[12] , \u_black_pixel_avg/black_pixel_count[13] , 
        \u_black_pixel_avg/black_pixel_count[14] , \u_black_pixel_avg/black_pixel_count[15] , 
        \u_black_pixel_avg/black_pixel_count[16] , \u_black_pixel_avg/black_pixel_count[17] , 
        \u_black_pixel_avg/black_pixel_count[18] , \u_black_pixel_avg/black_pixel_count[19] , 
        \u_black_pixel_avg/black_pixel_count[20] , \u_black_pixel_avg/black_pixel_count[21] , 
        \u_black_pixel_avg/black_pixel_count[22] , \u_black_pixel_avg/black_pixel_count[23] , 
        \u_black_pixel_avg/black_pixel_count[24] , \u_black_pixel_avg/black_pixel_count[25] , 
        \u_black_pixel_avg/black_pixel_count[26] , \u_black_pixel_avg/black_pixel_count[27] , 
        \u_black_pixel_avg/black_pixel_count[28] , \u_black_pixel_avg/black_pixel_count[29] , 
        \u_black_pixel_avg/black_pixel_count[30] , \u_black_pixel_avg/black_pixel_count[31] , 
        \x_avg_black[6] , \x_avg_black[7] , \x_avg_black[8] , \x_avg_black[9] , 
        \x_avg_black[10] , \x_avg_black[11] , n1812, n1813, n1814, 
        n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
        n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
        n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
        n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
        n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, 
        n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
        n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
        n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
        n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, 
        n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, 
        n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
        n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
        n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
        n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, 
        n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, 
        n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
        n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
        n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
        n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
        n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
        n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
        n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
        n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
        n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, 
        n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
        n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
        n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
        n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
        n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, 
        n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, 
        n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
        n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
        n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
        n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, 
        n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
        n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
        n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, 
        n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
        n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
        n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
        n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
        n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, 
        n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, 
        n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, 
        n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
        n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
        n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
        n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
        n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, 
        n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, 
        n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
        n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, 
        n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, 
        n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
        n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
        n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
        n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, 
        n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, 
        n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, 
        n2295, n2296, n2297, n2298, n2299, n2300, n2367, n2368, 
        n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, 
        n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, 
        n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
        n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
        n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
        n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, 
        n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, 
        n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
        n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
        n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, 
        n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, 
        n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, 
        n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
        n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
        n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, 
        n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, 
        n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, 
        n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
        n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
        n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, 
        n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, 
        n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
        n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
        n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, 
        n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, 
        n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, 
        n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, 
        n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
        n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
        n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, 
        n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, 
        n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, 
        n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
        n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, 
        n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
        n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, 
        n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, 
        n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, 
        n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, 
        n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
        n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
        n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, 
        n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
        n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
        n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
        n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
        n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
        n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, 
        n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, 
        n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
        n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
        n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, 
        n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
        n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, 
        n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
        n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
        n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, 
        n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
        n2833, n2834, n2835, n2836, n2837, n2838, n2842, n2843, 
        n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, 
        n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
        n2860, n2861, n2862, n2863, n2919, n2920, n2921, n2922, 
        n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
        n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
        n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
        n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, 
        n3008, n3009, n3052, n3053, n3054, n3055, n3056, n3057, 
        n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, 
        n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
        n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
        n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
        n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
        n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, 
        n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
        n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
        n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
        n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, 
        n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, 
        n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
        n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
        n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
        n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, 
        n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, 
        n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
        n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
        n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
        n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, 
        n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, 
        n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
        n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, 
        n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
        n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, 
        n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, 
        n3276, n3277, n3278, n3287, n3288, n3289, n3290, n3291, 
        n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, 
        n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, 
        n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, 
        n3316, n3317, n3318, n3319, n3320, n3327, n3328, n3329, 
        n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, 
        n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, 
        n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
        \y_avg_black[3] , \y_avg_black[4] , \y_avg_black[5] , \y_avg_black[6] , 
        \y_avg_black[7] , \y_avg_black[8] , \y_avg_black[9] , \y_avg_black[10] , 
        \y_avg_black[11] , \u_black_pixel_avg/x_sum[2] , \u_black_pixel_avg/x_sum[3] , 
        \u_black_pixel_avg/x_sum[4] , \u_black_pixel_avg/x_sum[5] , \u_black_pixel_avg/x_sum[6] , 
        \u_black_pixel_avg/x_sum[7] , \u_black_pixel_avg/x_sum[8] , \u_black_pixel_avg/x_sum[9] , 
        \u_black_pixel_avg/x_sum[10] , \u_black_pixel_avg/x_sum[11] , \u_black_pixel_avg/x_sum[12] , 
        \u_black_pixel_avg/x_sum[13] , \u_black_pixel_avg/x_sum[14] , \u_black_pixel_avg/x_sum[15] , 
        \u_black_pixel_avg/x_sum[16] , \u_black_pixel_avg/x_sum[17] , \u_black_pixel_avg/x_sum[18] , 
        \u_black_pixel_avg/x_sum[19] , \u_black_pixel_avg/x_sum[20] , \u_black_pixel_avg/x_sum[21] , 
        \u_black_pixel_avg/x_sum[22] , \u_black_pixel_avg/x_sum[23] , \u_black_pixel_avg/x_sum[24] , 
        \u_black_pixel_avg/x_sum[25] , \u_black_pixel_avg/x_sum[26] , \u_black_pixel_avg/x_sum[27] , 
        \u_black_pixel_avg/x_sum[28] , \u_black_pixel_avg/x_sum[29] , \u_black_pixel_avg/x_sum[30] , 
        \u_black_pixel_avg/x_sum[31] , n3395, n3396, n3397, n3398, 
        n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
        n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, 
        n3415, \u_state_machine/key0_last , \u_state_machine/current_state.WAITING , 
        \u_state_machine/current_state.WORKING , \u_state_machine/counter_10s[0] , 
        \u_state_machine/key0_debounced , \u_state_machine/counter_10s[1] , 
        \u_state_machine/counter_10s[2] , \u_state_machine/counter_10s[3] , 
        \u_state_machine/counter_10s[4] , \u_state_machine/counter_10s[5] , 
        \u_state_machine/counter_10s[6] , \u_state_machine/counter_10s[7] , 
        \u_state_machine/counter_10s[8] , \u_state_machine/counter_10s[9] , 
        \u_state_machine/counter_10s[10] , \u_state_machine/counter_10s[11] , 
        \u_state_machine/counter_10s[12] , \u_state_machine/counter_10s[13] , 
        \u_state_machine/counter_10s[14] , \u_state_machine/counter_10s[15] , 
        \u_state_machine/counter_10s[16] , \u_state_machine/counter_10s[17] , 
        \u_state_machine/counter_10s[18] , \u_state_machine/counter_10s[19] , 
        \u_state_machine/counter_10s[20] , \u_state_machine/counter_10s[21] , 
        \u_state_machine/counter_10s[22] , \u_state_machine/counter_10s[23] , 
        \u_state_machine/counter_10s[24] , \u_state_machine/counter_10s[25] , 
        \u_state_machine/counter_10s[26] , n3464, n3465, \w_hdmi_txd0[0] , 
        \u_rgb2dvi/enc_0/acc[0] , n3468, n3469, \w_hdmi_txd0[4] , \w_hdmi_txd0[8] , 
        \w_hdmi_txd0[9] , \u_rgb2dvi/enc_0/acc[1] , \u_rgb2dvi/enc_0/acc[2] , 
        \u_rgb2dvi/enc_0/acc[3] , \u_rgb2dvi/enc_0/acc[4] , n3478, n3479, 
        \w_hdmi_txd1[0] , \u_rgb2dvi/enc_1/acc[0] , \w_hdmi_txd1[4] , 
        \w_hdmi_txd1[8] , \w_hdmi_txd1[9] , \u_rgb2dvi/enc_1/acc[1] , 
        \u_rgb2dvi/enc_1/acc[2] , \u_rgb2dvi/enc_1/acc[3] , \u_rgb2dvi/enc_1/acc[4] , 
        n3490, n3491, n3492, n3493, \w_hdmi_txd2[0] , \u_rgb2dvi/enc_2/acc[0] , 
        \w_hdmi_txd2[4] , \w_hdmi_txd2[9] , \u_rgb2dvi/enc_2/acc[1] , 
        \u_rgb2dvi/enc_2/acc[2] , \u_rgb2dvi/enc_2/acc[3] , \u_rgb2dvi/enc_2/acc[4] , 
        \r_hdmi_tx0_o[6] , \r_hdmi_tx0_o[7] , \r_hdmi_tx0_o[8] , \r_hdmi_tx0_o[9] , 
        \r_hdmi_tx1_o[6] , \r_hdmi_tx1_o[7] , \r_hdmi_tx1_o[8] , \r_hdmi_tx1_o[9] , 
        \r_hdmi_tx2_o[6] , \r_hdmi_tx2_o[7] , \r_hdmi_tx2_o[9] , \PowerOnResetCnt[1] , 
        \PowerOnResetCnt[2] , \PowerOnResetCnt[3] , \PowerOnResetCnt[4] , 
        \PowerOnResetCnt[5] , \PowerOnResetCnt[6] , \PowerOnResetCnt[7] , 
        n642, n643, n644, n12160, n647, n648, n649, n650, n651, 
        n652, n653, n654, n3818, n3819, n3820, n3821, n3822, 
        n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, 
        n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, 
        n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, 
        n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, 
        n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
        n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, 
        n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, 
        n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, 
        n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, 
        n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, 
        n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, 
        n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
        n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, 
        n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, 
        n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, 
        n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, 
        n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, 
        n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, 
        n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, 
        n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, 
        n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, 
        n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, 
        n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, 
        n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, 
        n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, 
        n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, 
        n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
        n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, 
        n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, 
        n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, 
        n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, 
        n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
        n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, 
        n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, 
        n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, 
        n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, 
        n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
        n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
        n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, 
        n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, 
        n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, 
        n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
        n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, 
        n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, 
        n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
        n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, 
        n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
        n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, 
        n4207, n4208, n4209, n4210, n4211, n4212, n4220, n4221, 
        n4222, n4224, n4226, n4228, n4230, n4232, n4234, n4235, 
        n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, 
        n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, 
        n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, 
        n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
        n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, 
        n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
        n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, 
        n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, 
        n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
        n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, 
        n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
        n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, 
        n4332, n4333, n4334, n4335, n4349, n4350, n4351, n4352, 
        n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, 
        n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, 
        n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, 
        n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
        n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, 
        n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, 
        n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
        n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, 
        n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, 
        n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, 
        n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
        n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, 
        n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, 
        n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, 
        n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, 
        n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, 
        n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
        n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, 
        n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, 
        n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
        n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, 
        n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, 
        n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, 
        n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, 
        n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, 
        n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, 
        n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, 
        n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, 
        n4577, n4578, n4579, n4580, n4581, n4582, \Axi0ResetReg[1] , 
        \Axi0ResetReg[0] , \reduce_nand_9/n7 , DdrInitDone, w_XYCrop0_frame_vsync, 
        \w_XYCrop0_frame_Gray[0] , w_XYCrop0_frame_href, w_XYCrop0_frame_de, 
        \ResetShiftReg[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/n58 , \U0_DDR_Reset/u_ddr_reset_sequencer/n89 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/n92 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] , \U0_DDR_Reset/u_ddr_reset_sequencer/n57 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n91 , \U0_DDR_Reset/u_ddr_reset_sequencer/n56 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n55 , \U0_DDR_Reset/u_ddr_reset_sequencer/n54 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n53 , \U0_DDR_Reset/u_ddr_reset_sequencer/n52 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n51 , \U0_DDR_Reset/u_ddr_reset_sequencer/n50 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n49 , \U0_DDR_Reset/u_ddr_reset_sequencer/n48 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n47 , \U0_DDR_Reset/u_ddr_reset_sequencer/n46 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n45 , \U0_DDR_Reset/u_ddr_reset_sequencer/n44 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n43 , \U0_DDR_Reset/u_ddr_reset_sequencer/n42 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n41 , \U0_DDR_Reset/u_ddr_reset_sequencer/n40 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n39 , \U0_DDR_Reset/u_ddr_reset_sequencer/n38 , 
        \u_i2c_timing_ctrl_16bit/n158 , \u_i2c_timing_ctrl_16bit/n189 , 
        \u_i2c_timing_ctrl_16bit/n159 , \u_i2c_timing_ctrl_16bit/n160 , 
        \u_i2c_timing_ctrl_16bit/n241 , \u_i2c_timing_ctrl_16bit/n374 , 
        \u_i2c_timing_ctrl_16bit/n383 , \u_i2c_timing_ctrl_16bit/n63 , \u_i2c_timing_ctrl_16bit/n64 , 
        \u_i2c_timing_ctrl_16bit/n369 , \u_i2c_timing_ctrl_16bit/n157 , 
        \u_i2c_timing_ctrl_16bit/n156 , \u_i2c_timing_ctrl_16bit/n155 , 
        \u_i2c_timing_ctrl_16bit/n154 , \u_i2c_timing_ctrl_16bit/n153 , 
        \u_i2c_timing_ctrl_16bit/n152 , \u_i2c_timing_ctrl_16bit/n151 , 
        \u_i2c_timing_ctrl_16bit/n150 , \u_i2c_timing_ctrl_16bit/n149 , 
        \u_i2c_timing_ctrl_16bit/n148 , \u_i2c_timing_ctrl_16bit/n147 , 
        \u_i2c_timing_ctrl_16bit/n146 , \u_i2c_timing_ctrl_16bit/n145 , 
        \u_i2c_timing_ctrl_16bit/n144 , \u_i2c_timing_ctrl_16bit/n143 , 
        \u_i2c_timing_ctrl_16bit/n188 , \u_i2c_timing_ctrl_16bit/n187 , 
        \u_i2c_timing_ctrl_16bit/n186 , \u_i2c_timing_ctrl_16bit/n240 , 
        \u_i2c_timing_ctrl_16bit/n239 , \u_i2c_timing_ctrl_16bit/n238 , 
        \u_i2c_timing_ctrl_16bit/n237 , \u_i2c_timing_ctrl_16bit/n236 , 
        \u_i2c_timing_ctrl_16bit/n235 , \u_i2c_timing_ctrl_16bit/n234 , 
        \u_i2c_timing_ctrl_16bit/n233 , \u_i2c_timing_ctrl_16bit/n373 , 
        \u_i2c_timing_ctrl_16bit/n372 , \u_i2c_timing_ctrl_16bit/n371 , 
        \u_i2c_timing_ctrl_16bit/n382 , \u_i2c_timing_ctrl_16bit/n381 , 
        \u_i2c_timing_ctrl_16bit/n380 , \u_i2c_timing_ctrl_16bit/n379 , 
        \u_i2c_timing_ctrl_16bit/n378 , \u_i2c_timing_ctrl_16bit/n377 , 
        \u_i2c_timing_ctrl_16bit/n376 , \u_i2c_timing_ctrl_16bit/n62 , \u_i2c_timing_ctrl_16bit/n61 , 
        \u_i2c_timing_ctrl_16bit/n60 , \u_i2c_timing_ctrl_16bit/n59 , \u_i2c_timing_ctrl_16bit/n58 , 
        \u_i2c_timing_ctrl_16bit/n57 , \u_i2c_timing_ctrl_16bit/n56 , \u_i2c_timing_ctrl_16bit/n55 , 
        \u_i2c_timing_ctrl_16bit/n54 , \u_i2c_timing_ctrl_16bit/n53 , \u_i2c_timing_ctrl_16bit/n52 , 
        \u_i2c_timing_ctrl_16bit/n51 , \u_i2c_timing_ctrl_16bit/n50 , \u_i2c_timing_ctrl_16bit/n49 , 
        \u_i2c_timing_ctrl_16bit/n48 , \u_i2c_timing_ctrl_16bit/n47 , \u_i2c_timing_ctrl_16bit/n46 , 
        \u_i2c_timing_ctrl_16bit/n45 , \u_i2c_timing_ctrl_16bit/n44 , \u_i2c_timing_ctrl_16bit/n43 , 
        \u_i2c_timing_ctrl_16bit/n42 , \u_i2c_timing_ctrl_16bit/n41 , \u_i2c_timing_ctrl_16bit/n40 , 
        \u_i2c_timing_ctrl_16bit/n39 , \u_i2c_timing_ctrl_16bit/n38 , \u_Sensor_Image_XYCrop_0/n42 , 
        \u_Sensor_Image_XYCrop_0/n43 , \u_Sensor_Image_XYCrop_0/n44 , \u_Sensor_Image_XYCrop_0/n53 , 
        \u_Sensor_Image_XYCrop_0/n45 , \u_Sensor_Image_XYCrop_0/n46 , \u_Sensor_Image_XYCrop_0/n47 , 
        \u_Sensor_Image_XYCrop_0/n48 , \u_Sensor_Image_XYCrop_0/n49 , \u_Sensor_Image_XYCrop_0/n50 , 
        \u_Sensor_Image_XYCrop_0/n51 , \u_Sensor_Image_XYCrop_0/w_image_out_href , 
        \u_Sensor_Image_XYCrop_0/n52 , \axi4_awar_mux/n50 , \axi4_awar_mux/n131 , 
        \axi4_awar_mux/n52 , \axi4_awar_mux/n55 , \axi4_awar_mux/n49 , 
        \u_axi4_ctrl_0/n119 , \u_axi4_ctrl_0/n116 , \u_axi4_ctrl_0/n117 , 
        \u_axi4_ctrl_0/n120 , \u_axi4_ctrl_0/n265 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int , \u_axi4_ctrl_0/n290 , 
        \u_axi4_ctrl_0/n291 , \u_axi4_ctrl_0/n258 , \u_axi4_ctrl_0/n260 , 
        \u_axi4_ctrl_0/n346 , \u_axi4_ctrl_0/n267 , \u_axi4_ctrl_0/n266 , 
        \u_axi4_ctrl_0/n2649 , \u_axi4_ctrl_0/r_w_rst , lcd_vs, \u_axi4_ctrl_0/n1074 , 
        \u_axi4_ctrl_0/n2551 , \u_axi4_ctrl_0/n1075 , \u_axi4_ctrl_0/equal_138/n9 , 
        \u_axi4_ctrl_0/w_rfifo_rst , \u_axi4_ctrl_0/n2670 , \u_axi4_ctrl_0/r_rfifo_rst_rclk , 
        \u_axi4_ctrl_0/equal_160/n3 , \u_axi4_ctrl_0/n1730 , \u_axi4_ctrl_0/select_190/Select_1/n3 , 
        \u_axi4_ctrl_0/n1732 , \u_axi4_ctrl_0/n1733 , \u_axi4_ctrl_0/n1734 , 
        \u_axi4_ctrl_0/equal_189/n5 , \u_axi4_ctrl_0/n264 , \u_axi4_ctrl_0/n2777 , 
        \u_axi4_ctrl_0/n256 , \u_axi4_ctrl_0/n289 , \u_axi4_ctrl_0/n288 , 
        \u_axi4_ctrl_0/n287 , \u_axi4_ctrl_0/n286 , \u_axi4_ctrl_0/n285 , 
        \u_axi4_ctrl_0/n284 , \u_axi4_ctrl_0/n283 , \u_axi4_ctrl_0/n282 , 
        \u_axi4_ctrl_0/n281 , \u_axi4_ctrl_0/n280 , \u_axi4_ctrl_0/n279 , 
        \u_axi4_ctrl_0/n278 , \u_axi4_ctrl_0/n277 , \u_axi4_ctrl_0/n276 , 
        \u_axi4_ctrl_0/n275 , \u_axi4_ctrl_0/n274 , \u_axi4_ctrl_0/n273 , 
        \u_axi4_ctrl_0/n272 , \u_axi4_ctrl_0/n271 , \u_axi4_ctrl_0/n270 , 
        \u_axi4_ctrl_0/n269 , \u_axi4_ctrl_0/n345 , \u_axi4_ctrl_0/n344 , 
        \u_axi4_ctrl_0/n343 , \u_axi4_ctrl_0/n342 , \u_axi4_ctrl_0/n341 , 
        \u_axi4_ctrl_0/n340 , \u_axi4_ctrl_0/n339 , \u_axi4_ctrl_0/n766 , 
        \u_axi4_ctrl_0/n765 , \u_axi4_ctrl_0/n764 , \u_axi4_ctrl_0/n763 , 
        \u_axi4_ctrl_0/n762 , \u_axi4_ctrl_0/n761 , \u_axi4_ctrl_0/n760 , 
        \u_axi4_ctrl_0/n759 , \u_axi4_ctrl_0/n758 , \u_axi4_ctrl_0/n757 , 
        \u_axi4_ctrl_0/n756 , \u_axi4_ctrl_0/n755 , \u_axi4_ctrl_0/n754 , 
        \u_axi4_ctrl_0/n753 , \u_axi4_ctrl_0/n752 , \u_axi4_ctrl_0/n751 , 
        \u_axi4_ctrl_0/n750 , \u_axi4_ctrl_0/n749 , \u_axi4_ctrl_0/n748 , 
        \u_axi4_ctrl_0/n747 , \u_axi4_ctrl_0/n746 , \u_axi4_ctrl_0/n745 , 
        \u_axi4_ctrl_0/n744 , \u_axi4_ctrl_0/n743 , \u_axi4_ctrl_0/n742 , 
        \u_axi4_ctrl_0/n741 , \u_axi4_ctrl_0/n740 , \u_axi4_ctrl_0/n739 , 
        \u_axi4_ctrl_0/n738 , \u_axi4_ctrl_0/n737 , \u_axi4_ctrl_0/n736 , 
        \u_axi4_ctrl_0/n735 , \u_axi4_ctrl_0/n734 , \u_axi4_ctrl_0/n733 , 
        \u_axi4_ctrl_0/n732 , \u_axi4_ctrl_0/n731 , \u_axi4_ctrl_0/n730 , 
        \u_axi4_ctrl_0/n729 , \u_axi4_ctrl_0/n728 , \u_axi4_ctrl_0/n727 , 
        \u_axi4_ctrl_0/n726 , \u_axi4_ctrl_0/n725 , \u_axi4_ctrl_0/n724 , 
        \u_axi4_ctrl_0/n723 , \u_axi4_ctrl_0/n722 , \u_axi4_ctrl_0/n721 , 
        \u_axi4_ctrl_0/n720 , \u_axi4_ctrl_0/n719 , \u_axi4_ctrl_0/n718 , 
        \u_axi4_ctrl_0/n717 , \u_axi4_ctrl_0/n716 , \u_axi4_ctrl_0/n715 , 
        \u_axi4_ctrl_0/n714 , \u_axi4_ctrl_0/n713 , \u_axi4_ctrl_0/n712 , 
        \u_axi4_ctrl_0/n711 , \u_axi4_ctrl_0/n710 , \u_axi4_ctrl_0/n709 , 
        \u_axi4_ctrl_0/n708 , \u_axi4_ctrl_0/n707 , \u_axi4_ctrl_0/n706 , 
        \u_axi4_ctrl_0/n705 , \u_axi4_ctrl_0/n704 , \u_axi4_ctrl_0/n703 , 
        \u_axi4_ctrl_0/n702 , \u_axi4_ctrl_0/n701 , \u_axi4_ctrl_0/n700 , 
        \u_axi4_ctrl_0/n699 , \u_axi4_ctrl_0/n698 , \u_axi4_ctrl_0/n697 , 
        \u_axi4_ctrl_0/n696 , \u_axi4_ctrl_0/n695 , \u_axi4_ctrl_0/n694 , 
        \u_axi4_ctrl_0/n693 , \u_axi4_ctrl_0/n692 , \u_axi4_ctrl_0/n691 , 
        \u_axi4_ctrl_0/n690 , \u_axi4_ctrl_0/n689 , \u_axi4_ctrl_0/n688 , 
        \u_axi4_ctrl_0/n687 , \u_axi4_ctrl_0/n686 , \u_axi4_ctrl_0/n685 , 
        \u_axi4_ctrl_0/n684 , \u_axi4_ctrl_0/n683 , \u_axi4_ctrl_0/n682 , 
        \u_axi4_ctrl_0/n681 , \u_axi4_ctrl_0/n680 , \u_axi4_ctrl_0/n679 , 
        \u_axi4_ctrl_0/n678 , \u_axi4_ctrl_0/n677 , \u_axi4_ctrl_0/n676 , 
        \u_axi4_ctrl_0/n675 , \u_axi4_ctrl_0/n674 , \u_axi4_ctrl_0/n673 , 
        \u_axi4_ctrl_0/n672 , \u_axi4_ctrl_0/n671 , \u_axi4_ctrl_0/n670 , 
        \u_axi4_ctrl_0/n669 , \u_axi4_ctrl_0/n668 , \u_axi4_ctrl_0/n667 , 
        \u_axi4_ctrl_0/n666 , \u_axi4_ctrl_0/n665 , \u_axi4_ctrl_0/n664 , 
        \u_axi4_ctrl_0/n663 , \u_axi4_ctrl_0/n662 , \u_axi4_ctrl_0/n661 , 
        \u_axi4_ctrl_0/n660 , \u_axi4_ctrl_0/n659 , \u_axi4_ctrl_0/n658 , 
        \u_axi4_ctrl_0/n657 , \u_axi4_ctrl_0/n656 , \u_axi4_ctrl_0/n655 , 
        \u_axi4_ctrl_0/n654 , \u_axi4_ctrl_0/n653 , \u_axi4_ctrl_0/n652 , 
        \u_axi4_ctrl_0/n651 , \u_axi4_ctrl_0/n650 , \u_axi4_ctrl_0/n649 , 
        \u_axi4_ctrl_0/n648 , \u_axi4_ctrl_0/n647 , \u_axi4_ctrl_0/n2656 , 
        \u_axi4_ctrl_0/n2661 , \u_axi4_ctrl_0/n2666 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n71 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n152 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n184 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n194 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n151 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n150 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n149 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n148 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n147 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n146 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n145 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n144 , 
        n5390, \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n183 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n182 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n181 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n180 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n179 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n178 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n177 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n176 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n193 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n192 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n191 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n190 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n189 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n188 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n187 , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n186 , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl_0/n1073 , \u_axi4_ctrl_0/n1072 , \u_axi4_ctrl_0/n1071 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n71 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n152 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n184 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n194 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n151 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n150 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n149 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n148 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n147 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n146 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n145 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n144 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n183 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n182 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n181 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n180 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n179 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n178 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n177 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n176 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n193 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n192 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n191 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n190 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n189 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n188 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n187 , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n186 , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl_0/n2677 , \u_axi4_ctrl_0/n2682 , \u_axi4_ctrl_0/n1507 , 
        \u_axi4_ctrl_0/n1506 , \u_axi4_ctrl_0/n1505 , \u_axi4_ctrl_0/n1504 , 
        \u_axi4_ctrl_0/n1503 , \u_axi4_ctrl_0/n1502 , \u_axi4_ctrl_0/n1501 , 
        \u_axi4_ctrl_0/n1500 , \u_axi4_ctrl_0/n1499 , \u_axi4_ctrl_0/n1498 , 
        \u_axi4_ctrl_0/n1497 , \u_axi4_ctrl_0/n1496 , \u_axi4_ctrl_0/n1495 , 
        \u_axi4_ctrl_0/n1494 , \u_axi4_ctrl_0/n1493 , \u_axi4_ctrl_0/n1492 , 
        \u_axi4_ctrl_0/n1491 , \u_axi4_ctrl_0/n1490 , \u_axi4_ctrl_0/n1489 , 
        \u_axi4_ctrl_0/n1488 , \u_axi4_ctrl_0/n1487 , \u_axi4_ctrl_0/n1486 , 
        \u_axi4_ctrl_0/n1485 , \u_axi4_ctrl_0/n1484 , \u_axi4_ctrl_0/n1483 , 
        \u_axi4_ctrl_0/n1482 , \u_axi4_ctrl_0/n1481 , \u_axi4_ctrl_0/n1480 , 
        \u_axi4_ctrl_0/n1479 , \u_axi4_ctrl_0/n1478 , \u_axi4_ctrl_0/n1477 , 
        \u_axi4_ctrl_0/n1476 , \u_axi4_ctrl_0/n1475 , \u_axi4_ctrl_0/n1474 , 
        \u_axi4_ctrl_0/n1473 , \u_axi4_ctrl_0/n1472 , \u_axi4_ctrl_0/n1471 , 
        \u_axi4_ctrl_0/n1470 , \u_axi4_ctrl_0/n1469 , \u_axi4_ctrl_0/n1468 , 
        \u_axi4_ctrl_0/n1467 , \u_axi4_ctrl_0/n1466 , \u_axi4_ctrl_0/n1465 , 
        \u_axi4_ctrl_0/n1464 , \u_axi4_ctrl_0/n1463 , \u_axi4_ctrl_0/n1462 , 
        \u_axi4_ctrl_0/n1461 , \u_axi4_ctrl_0/n1460 , \u_axi4_ctrl_0/n1459 , 
        \u_axi4_ctrl_0/n1458 , \u_axi4_ctrl_0/n1457 , \u_axi4_ctrl_0/n1456 , 
        \u_axi4_ctrl_0/n1455 , \u_axi4_ctrl_0/n1454 , \u_axi4_ctrl_0/n1453 , 
        \u_axi4_ctrl_0/n1452 , \u_axi4_ctrl_0/n1451 , \u_axi4_ctrl_0/n1450 , 
        \u_axi4_ctrl_0/n1449 , \u_axi4_ctrl_0/n1448 , \u_axi4_ctrl_0/n1447 , 
        \u_axi4_ctrl_0/n1446 , \u_axi4_ctrl_0/n1445 , \u_axi4_ctrl_0/n1444 , 
        \u_axi4_ctrl_0/n1443 , \u_axi4_ctrl_0/n1442 , \u_axi4_ctrl_0/n1441 , 
        \u_axi4_ctrl_0/n1440 , \u_axi4_ctrl_0/n1439 , \u_axi4_ctrl_0/n1438 , 
        \u_axi4_ctrl_0/n1437 , \u_axi4_ctrl_0/n1436 , \u_axi4_ctrl_0/n1435 , 
        \u_axi4_ctrl_0/n1434 , \u_axi4_ctrl_0/n1433 , \u_axi4_ctrl_0/n1432 , 
        \u_axi4_ctrl_0/n1431 , \u_axi4_ctrl_0/n1430 , \u_axi4_ctrl_0/n1429 , 
        \u_axi4_ctrl_0/n1428 , \u_axi4_ctrl_0/n1427 , \u_axi4_ctrl_0/n1426 , 
        \u_axi4_ctrl_0/n1425 , \u_axi4_ctrl_0/n1424 , \u_axi4_ctrl_0/n1423 , 
        \u_axi4_ctrl_0/n1422 , \u_axi4_ctrl_0/n1421 , \u_axi4_ctrl_0/n1420 , 
        \u_axi4_ctrl_0/n1419 , \u_axi4_ctrl_0/n1418 , \u_axi4_ctrl_0/n1417 , 
        \u_axi4_ctrl_0/n1416 , \u_axi4_ctrl_0/n1415 , \u_axi4_ctrl_0/n1414 , 
        \u_axi4_ctrl_0/n1413 , \u_axi4_ctrl_0/n1412 , \u_axi4_ctrl_0/n1411 , 
        \u_axi4_ctrl_0/n1410 , \u_axi4_ctrl_0/n1409 , \u_axi4_ctrl_0/n1408 , 
        \u_axi4_ctrl_0/n1407 , \u_axi4_ctrl_0/n1406 , \u_axi4_ctrl_0/n1405 , 
        \u_axi4_ctrl_0/n1404 , \u_axi4_ctrl_0/n1403 , \u_axi4_ctrl_0/n1402 , 
        \u_axi4_ctrl_0/n1401 , \u_axi4_ctrl_0/n1400 , \u_axi4_ctrl_0/n1399 , 
        \u_axi4_ctrl_0/n1398 , \u_axi4_ctrl_0/n1397 , \u_axi4_ctrl_0/n1396 , 
        \u_axi4_ctrl_0/n1395 , \u_axi4_ctrl_0/n1394 , \u_axi4_ctrl_0/n1393 , 
        \u_axi4_ctrl_0/n1392 , \u_axi4_ctrl_0/n1391 , \u_axi4_ctrl_0/n1390 , 
        \u_axi4_ctrl_0/n1389 , \u_axi4_ctrl_0/n1388 , \u_axi4_ctrl_0/n1387 , 
        \u_axi4_ctrl_0/n1386 , \u_axi4_ctrl_0/n1385 , \u_axi4_ctrl_0/n1384 , 
        \u_axi4_ctrl_0/n1383 , \u_axi4_ctrl_0/n1382 , \u_axi4_ctrl_0/n1381 , 
        \u_axi4_ctrl_0/n1380 , \u_lcd_driver/hcnt[0] , \u_axi4_ctrl_0/n1774 , 
        \u_axi4_ctrl_0/n1773 , \u_axi4_ctrl_0/n1772 , \u_axi4_ctrl_0/n1771 , 
        \u_axi4_ctrl_0/n1770 , \u_axi4_ctrl_0/n1769 , \u_axi4_ctrl_0/n1768 , 
        \u_axi4_ctrl_0/n1767 , \u_axi4_ctrl_0/n1766 , \u_axi4_ctrl_0/n1765 , 
        \u_axi4_ctrl_0/n1764 , \u_axi4_ctrl_0/n1763 , \u_axi4_ctrl_0/n1762 , 
        \u_axi4_ctrl_0/n1761 , \u_axi4_ctrl_0/n2772 , \u_lcd_driver/n96 , 
        \u_lcd_driver/n51 , \u_lcd_driver/n113 , \u_lcd_driver/n125 , 
        \u_lcd_driver/n194 , \u_lcd_driver/n34 , \u_lcd_driver/n95 , \u_lcd_driver/n94 , 
        \u_lcd_driver/n93 , \u_lcd_driver/n92 , \u_lcd_driver/n91 , \u_lcd_driver/n90 , 
        \u_lcd_driver/n89 , \u_lcd_driver/n88 , \u_lcd_driver/n87 , \u_lcd_driver/n86 , 
        \u_lcd_driver/n85 , n733, \u_lcd_driver/n33 , \u_lcd_driver/n32 , 
        \u_lcd_driver/n31 , \u_lcd_driver/n30 , \u_lcd_driver/n29 , \u_lcd_driver/n28 , 
        \u_lcd_driver/n27 , \u_lcd_driver/n26 , \u_lcd_driver/n25 , \u_lcd_driver/n24 , 
        \u_lcd_driver/n23 , \u_black_pixel_avg/n175 , \u_black_pixel_avg/n208 , 
        \u_black_pixel_avg/n141 , \u_black_pixel_avg/n142 , \u_black_pixel_avg/n174 , 
        \u_black_pixel_avg/n173 , \u_black_pixel_avg/n172 , \u_black_pixel_avg/n171 , 
        \u_black_pixel_avg/n170 , \u_black_pixel_avg/n169 , \u_black_pixel_avg/n168 , 
        \u_black_pixel_avg/n167 , \u_black_pixel_avg/n166 , \u_black_pixel_avg/n165 , 
        \u_black_pixel_avg/n164 , \u_black_pixel_avg/n163 , \u_black_pixel_avg/n162 , 
        \u_black_pixel_avg/n161 , \u_black_pixel_avg/n160 , \u_black_pixel_avg/n159 , 
        \u_black_pixel_avg/n158 , \u_black_pixel_avg/n157 , \u_black_pixel_avg/n156 , 
        \u_black_pixel_avg/n155 , \u_black_pixel_avg/n154 , \u_black_pixel_avg/n153 , 
        \u_black_pixel_avg/n152 , \u_black_pixel_avg/n151 , \u_black_pixel_avg/n150 , 
        \u_black_pixel_avg/n149 , \u_black_pixel_avg/n148 , \u_black_pixel_avg/n147 , 
        \u_black_pixel_avg/n146 , \u_black_pixel_avg/n145 , \u_black_pixel_avg/n144 , 
        \u_black_pixel_avg/n207 , \u_black_pixel_avg/n206 , \u_black_pixel_avg/n205 , 
        \u_black_pixel_avg/n204 , \u_black_pixel_avg/n203 , \u_black_pixel_avg/n202 , 
        \u_black_pixel_avg/n201 , \u_black_pixel_avg/n200 , \u_black_pixel_avg/n199 , 
        \u_black_pixel_avg/n198 , \u_black_pixel_avg/n197 , \u_black_pixel_avg/n196 , 
        \u_black_pixel_avg/n195 , \u_black_pixel_avg/n194 , \u_black_pixel_avg/n193 , 
        \u_black_pixel_avg/n192 , \u_black_pixel_avg/n191 , \u_black_pixel_avg/n190 , 
        \u_black_pixel_avg/n189 , \u_black_pixel_avg/n188 , \u_black_pixel_avg/n187 , 
        \u_black_pixel_avg/n186 , \u_black_pixel_avg/n185 , \u_black_pixel_avg/n184 , 
        \u_black_pixel_avg/n183 , \u_black_pixel_avg/n182 , \u_black_pixel_avg/n181 , 
        \u_black_pixel_avg/n180 , \u_black_pixel_avg/n179 , \u_black_pixel_avg/n178 , 
        \u_black_pixel_avg/n177 , \u_black_pixel_avg/n483 , \u_black_pixel_avg/n482 , 
        \u_black_pixel_avg/n481 , \u_black_pixel_avg/n480 , \u_black_pixel_avg/n479 , 
        \u_black_pixel_avg/n478 , n6202, n6206, n6209, n6212, n6215, 
        n6217, n6220, n6223, n6225, n6227, n6230, n6233, n6235, 
        n6237, n6239, n6242, n6245, n6247, n6249, n6251, n6253, 
        n6256, n6259, n6261, n6263, n6265, n6267, n6269, n6272, 
        n6275, n6277, n6279, n6281, n6283, n6285, n6287, n6290, 
        n6293, n6295, n6297, n6299, n6301, n6303, n6305, n6307, 
        n6310, n6313, n6315, n6317, n6319, n6321, n6323, n6325, 
        n6327, n6329, n6332, n6335, n6337, n6339, n6341, n6343, 
        n6345, n6347, n6349, n6351, n6353, n6356, n6359, n6361, 
        n6363, n6365, n6367, n6369, n6371, n6373, n6375, n6377, 
        n6379, n6382, n6385, n6387, n6389, n6391, n6393, n6395, 
        n6397, n6399, n6401, n6403, n6405, n6407, n6410, n6413, 
        n6415, n6417, n6419, n6421, n6423, n6425, n6427, n6429, 
        n6431, n6433, n6435, n6437, n6440, n6443, n6445, n6447, 
        n6449, n6451, n6453, n6455, n6457, n6459, n6461, n6463, 
        n6465, n6467, n6469, n6472, n6475, n6477, n6479, n6481, 
        n6483, n6485, n6487, n6489, n6491, n6493, n6495, n6497, 
        n6499, n6501, n6503, n6506, n6508, n6510, n6512, n6514, 
        n6516, n6518, n6520, n6522, n6524, n6526, n6528, n6530, 
        n6532, n6534, n6537, n6539, n6541, n6543, n6545, n6547, 
        n6549, n6551, n6553, n6555, n6557, n6559, n6561, n6563, 
        n6566, n6568, n6570, n6572, n6574, n6576, n6578, n6580, 
        n6582, n6584, n6586, n6588, n6590, n6593, n6595, n6597, 
        n6599, n6601, n6603, n6605, n6607, n6609, n6611, n6613, 
        n6615, n6618, n6620, n6622, n6624, n6626, n6628, n6630, 
        n6632, n6634, n6636, n6638, n6641, n6643, n6645, n6647, 
        n6649, n6651, n6653, n6655, n6657, n6659, n6662, n6664, 
        n6666, n6668, n6670, n6672, n6674, n6676, n6678, n6681, 
        n6683, n6685, n6687, n6689, n6691, n6693, n6695, n6698, 
        n6700, n6702, n6704, n6706, n6759, n6762, n6764, n6767, 
        n6769, n6771, n6774, n6776, n6778, n6780, n6783, n6785, 
        n6787, n6789, n6791, n6794, n6796, n6798, n6800, n6802, 
        n6804, n6807, n6809, n6811, n6813, n6815, n6817, n6819, 
        n6822, n6824, n6826, n6828, n6830, n6832, n6834, n6836, 
        n6839, n6841, n6843, n6845, n6847, n6849, n6851, n6853, 
        n6855, n6858, n6860, n6862, n6864, n6866, n6868, n6870, 
        n6872, n6874, n6876, n6879, n6881, n6883, n6885, n6887, 
        n6889, n6891, n6893, n6895, n6897, n6899, n6902, n6904, 
        n6906, n6908, n6910, n6912, n6914, n6916, n6918, n6920, 
        n6922, n6924, n6927, n6929, n6931, n6933, n6935, n6937, 
        n6939, n6941, n6943, n6945, n6947, n6949, n6951, n6954, 
        n6956, n6958, n6960, n6962, n6964, n6966, n6968, n6970, 
        n6972, n6974, n6976, n6978, n6980, n6983, n6985, n6987, 
        n6989, n6991, n6993, n6995, n6997, n6999, n7001, n7003, 
        n7005, n7007, n7009, n7011, n7014, n7016, n7018, n7020, 
        n7022, n7024, n7026, n7028, n7030, n7032, n7034, n7036, 
        n7038, n7040, n7042, n7044, n7047, n7049, n7051, n7053, 
        n7055, n7057, n7059, n7061, n7063, n7065, n7067, n7069, 
        n7071, n7073, n7075, n7078, n7080, n7082, n7084, n7086, 
        n7088, n7090, n7092, n7094, n7096, n7098, n7100, n7102, 
        n7104, n7107, n7109, n7111, n7113, n7115, n7117, n7119, 
        n7121, n7123, n7125, n7127, n7129, n7131, n7134, n7136, 
        n7138, n7140, n7142, n7144, n7146, n7148, n7150, n7152, 
        n7154, n7156, n7160, n7163, n7166, n7169, n7174, n7177, 
        n7180, n7183, n7185, n7187, n7189, n7191, n7193, n7195, 
        n7197, n7199, n7201, n7203, n7205, n7221, n7226, n7229, 
        n7232, n7235, n7245, n7247, n7249, n7251, n7253, n7255, 
        n7257, n7259, n7261, n7263, n7334, n7336, n7338, n7340, 
        n7342, n7344, n7346, n7348, n7350, n7401, n7403, n7405, 
        n7407, n7409, n7411, n7413, n7415, n7417, n7419, n7421, 
        n7424, n7426, n7428, n7430, n7432, n7434, n7436, n7438, 
        n7440, n7442, n7444, n7446, n7448, n7450, n7452, n7454, 
        n7456, n7458, n7460, n7464, n7466, n7468, n7470, n7472, 
        n7474, n7476, n7478, n7480, n7482, n7484, n7486, n7488, 
        n7491, n7493, n7495, n7497, n7499, n7501, n7503, n7505, 
        n7507, n7509, n7511, n7513, n7515, n7517, n7519, n7521, 
        n7523, n7525, n7527, n7529, n7531, n7533, n7535, n7537, 
        n7539, n7541, n7543, n7545, n7547, n7549, n7551, n7554, 
        n7556, n7558, n7560, n7562, n7564, n7566, n7568, n7570, 
        n7572, n7574, n7576, n7578, n7580, n7582, n7584, n7586, 
        n7588, n7590, n7592, n7594, n7596, n7598, n7600, n7602, 
        n7604, n7606, n7608, n7610, n7613, n7615, n7617, n7619, 
        n7621, n7623, n7625, n7627, n7629, n7631, n7633, n7635, 
        n7637, n7639, n7641, n7643, n7645, n7647, n7649, n7651, 
        n7653, n7655, n7666, n7668, n7670, n7672, n7674, n7676, 
        n7678, n7680, n7682, n7684, n7686, n7688, n7690, n7692, 
        n7701, n7703, n7705, n7707, n7709, n7711, n7713, n7715, 
        n7717, n7719, n7721, n7723, n7725, n7727, n7729, n7731, 
        n7733, n7735, n7742, n7744, n7746, n7748, n7750, n7752, 
        n7754, n7756, n7758, n7760, n7762, n7764, \u_black_pixel_avg/n499 , 
        \u_black_pixel_avg/n498 , \u_black_pixel_avg/n497 , \u_black_pixel_avg/n496 , 
        \u_black_pixel_avg/n495 , \u_black_pixel_avg/n494 , \u_black_pixel_avg/n493 , 
        \u_black_pixel_avg/n492 , \u_black_pixel_avg/n491 , \u_black_pixel_avg/n140 , 
        \u_black_pixel_avg/n139 , \u_black_pixel_avg/n138 , \u_black_pixel_avg/n137 , 
        \u_black_pixel_avg/n136 , \u_black_pixel_avg/n135 , \u_black_pixel_avg/n134 , 
        \u_black_pixel_avg/n133 , \u_black_pixel_avg/n132 , \u_black_pixel_avg/n131 , 
        \u_black_pixel_avg/n130 , \u_black_pixel_avg/n129 , \u_black_pixel_avg/n128 , 
        \u_black_pixel_avg/n127 , \u_black_pixel_avg/n126 , \u_black_pixel_avg/n125 , 
        \u_black_pixel_avg/n124 , \u_black_pixel_avg/n123 , \u_black_pixel_avg/n122 , 
        \u_black_pixel_avg/n121 , \u_black_pixel_avg/n120 , \u_black_pixel_avg/n119 , 
        \u_black_pixel_avg/n118 , \u_black_pixel_avg/n117 , \u_black_pixel_avg/n116 , 
        \u_black_pixel_avg/n115 , \u_black_pixel_avg/n114 , \u_black_pixel_avg/n113 , 
        \u_black_pixel_avg/n112 , \u_black_pixel_avg/n111 , n7811, n7813, 
        n7815, n7817, n7819, n7821, n7823, n7825, n7827, n7829, 
        n7831, n7833, \u_state_machine/next_state.WAITING , \u_state_machine/n113 , 
        \u_state_machine/next_state.WORKING , \u_state_machine/n99 , \u_state_machine/equal_19/n3 , 
        \u_state_machine/n114 , \u_state_machine/n115 , \u_state_machine/n116 , 
        \u_state_machine/n150 , \u_state_machine/n5 , \u_state_machine/n112 , 
        \u_state_machine/n111 , \u_state_machine/n110 , \u_state_machine/n109 , 
        \u_state_machine/n108 , \u_state_machine/n107 , \u_state_machine/n106 , 
        \u_state_machine/n98 , \u_state_machine/n97 , \u_state_machine/n96 , 
        \u_state_machine/n95 , \u_state_machine/n94 , \u_state_machine/n93 , 
        \u_state_machine/n92 , \u_state_machine/n91 , \u_state_machine/n90 , 
        \u_state_machine/n89 , \u_state_machine/n88 , \u_state_machine/n87 , 
        \u_state_machine/n86 , \u_state_machine/n85 , \u_state_machine/n84 , 
        \u_state_machine/n83 , \u_state_machine/n82 , \u_state_machine/n81 , 
        \u_state_machine/n80 , \u_state_machine/n79 , \u_state_machine/n78 , 
        \u_state_machine/n77 , \u_state_machine/n76 , \u_state_machine/n75 , 
        \u_state_machine/n74 , \u_state_machine/n73 , \u_rgb2dvi/enc_0/n869 , 
        \u_rgb2dvi/enc_0/n770 , \u_rgb2dvi/enc_0/n806 , \u_rgb2dvi/enc_0/n812 , 
        \u_rgb2dvi/enc_1/q_out[9] , \u_rgb2dvi/enc_2/q_out[9] , \r_hdmi_txc_o[9] , 
        n8196, n8198, n8200, n8202, n8204, n8206, n8208, n8210, 
        n8212, n8214, n8216, n8218, n8220, n8224, n8226, n8228, 
        n8230, n8232, n8234, n8236, n8238, n8240, n8242, n8244, 
        n8246, n8248, n8250, n8252, n8254, n8256, n8258, n8260, 
        n8262, n8264, n8266, n8268, n8270, n8272, n8274, n8276, 
        n8278, n8280, n8282, n8284, n8286, n8288, n8290, n8292, 
        n8294, n8296, n8298, n8300, n8302, n8304, n8306, n8308, 
        n8310, n8312, n8314, n8316, n8318, n8320, n8322, n8324, 
        n8326, n8328, n8330, n8332, n8334, n8336, n8338, n8340, 
        n8342, n8344, n8346, n8348, n8350, n8352, n8354, n8356, 
        n8358, n8360, n8362, n8364, n8366, n8368, n8370, n8372, 
        n8651, n8654, n8657, n8660, n8663, n8666, n8669, n8672, 
        \hdmi_clk1x_i~O , \Axi0Clk~O , \cmos_pclk~O , \hdmi_clk2x_i~O , 
        n12216, n12215, n12214, n12213, n12212, n12208, n12207, 
        n12206, n12205, n12204, n12203, n12202, n12201, n12200, 
        n12199, n12198, n12197, n12196, n12195, n12194, n12193, 
        n12192, n12191, n12190, n12189, n12188, n12187, n12186, 
        n12185, n12184, n12183, n12182, n12181, n12174, n12173, 
        n12172, n12171, n12170, n12169, n12168, n12167, n12166, 
        n12165, n12164, n12163, n12162, n12159, n12158, n12157, 
        n12156, n12155, n12154, n12153, n8971, n12152, n8974, 
        n12151, n12150, n12149, n12148, n12146, n12145, n12144, 
        n12143, n12142, n12141, n8988, n8989, n8990, n8991, n8992, 
        n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, 
        n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, 
        n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, 
        n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, 
        n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, 
        n9033, n9034, n9035, n9036, n9037, n9040, n9041, n9042, 
        n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, 
        n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, 
        n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, 
        n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, 
        n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, 
        n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, 
        n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, 
        n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, 
        n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, 
        n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, 
        n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, 
        n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9143, 
        n9145, n9149, n9150, n9151, n9152, n9153, n9154, n9155, 
        n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
        n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, 
        n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, 
        n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
        n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, 
        n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
        n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, 
        n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, 
        n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, 
        n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, 
        n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
        n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, 
        n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, 
        n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, 
        n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, 
        n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, 
        n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, 
        n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, 
        n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, 
        n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, 
        n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
        n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, 
        n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, 
        n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, 
        n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, 
        n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, 
        n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, 
        n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, 
        n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, 
        n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, 
        n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, 
        n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, 
        n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, 
        n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, 
        n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, 
        n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, 
        n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, 
        n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, 
        n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, 
        n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, 
        n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, 
        n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, 
        n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, 
        n9501, n9503, n9504, n9505, n9506, n9507, n9508, n9509, 
        n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, 
        n9518, n9519, n9520, n9523, n9524, n9525, n9526, n9527, 
        n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, 
        n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, 
        n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, 
        n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, 
        n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, 
        n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, 
        n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, 
        n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, 
        n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, 
        n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, 
        n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, 
        n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, 
        n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, 
        n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, 
        n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, 
        n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, 
        n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, 
        n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, 
        n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, 
        n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, 
        n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, 
        n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, 
        n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, 
        n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, 
        n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, 
        n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, 
        n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, 
        n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, 
        n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, 
        n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, 
        n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, 
        n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, 
        n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, 
        n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, 
        n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, 
        n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, 
        n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
        n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, 
        n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, 
        n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, 
        n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, 
        n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, 
        n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, 
        n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, 
        n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, 
        n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, 
        n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, 
        n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, 
        n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, 
        n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, 
        n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, 
        n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, 
        n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, 
        n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, 
        n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, 
        n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, 
        n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, 
        n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, 
        n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, 
        n10000, n10001, n10002, n10003, n10004, n10005, n10006, 
        n10007, n10008, n10009, n10010, n10011, n10012, n10013, 
        n10014, n10015, n10016, n10017, n10018, n10019, n10020, 
        n10021, n10022, n10023, n10024, n10025, n10026, n10027, 
        n10028, n10029, n10030, n10031, n10032, n10033, n10034, 
        n10035, n10036, n10037, n10038, n10039, n10040, n10041, 
        n10042, n10043, n10044, n10045, n10046, n10047, n10048, 
        n10049, n10050, n10051, n10052, n10053, n10054, n10055, 
        n10056, n10057, n10058, n10059, n10060, n10061, n10062, 
        n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
        n10070, n10071, n10072, n10073, n10074, n10075, n10076, 
        n10077, n10078, n10079, n10080, n10081, n10082, n10083, 
        n10084, n10085, n10086, n10087, n10088, n10089, n10090, 
        n10091, n10092, n10093, n10094, n10095, n10096, n10097, 
        n10098, n10099, n10100, n10101, n10102, n10103, n10104, 
        n10105, n10106, n10107, n10108, n10109, n10110, n10111, 
        n10112, n10113, n10114, n10115, n10116, n10117, n10118, 
        n10119, n10120, n10121, n10122, n10123, n10124, n10125, 
        n10126, n10127, n10128, n10129, n10130, n10131, n10132, 
        n10133, n10134, n10135, n10136, n10137, n10138, n10139, 
        n10140, n10141, n10142, n10143, n10144, n10145, n10146, 
        n10147, n10148, n10149, n10150, n10151, n10152, n10153, 
        n10154, n10155, n10156, n10157, n10158, n10159, n10160, 
        n10161, n10162, n10163, n10164, n10165, n10166, n10167, 
        n10168, n10169, n10170, n10171, n10172, n10173, n10174, 
        n10175, n10176, n10177, n10178, n10179, n10180, n10181, 
        n10182, n10183, n10184, n10185, n10186, n10187, n10188, 
        n10189, n10190, n10191, n10192, n10193, n10194, n10195, 
        n10196, n10197, n10198, n10199, n10200, n10201, n10202, 
        n10203, n10204, n10205, n10206, n10207, n10208, n10209, 
        n10210, n10211, n10212, n10213, n10214, n10215, n10216, 
        n10217, n10218, n10219, n10220, n10221, n10222, n10223, 
        n10224, n10225, n10226, n10227, n10228, n10229, n10230, 
        n10231, n10232, n10233, n10234, n10235, n10236, n10237, 
        n10238, n10239, n10240, n10241, n10242, n10243, n10244, 
        n10245, n10246, n10247, n10248, n10249, n10250, n10251, 
        n10252, n10253, n10254, n10255, n10256, n10257, n10258, 
        n10259, n10260, n10261, n10262, n10263, n10264, n10265, 
        n10266, n10267, n10268, n10269, n10270, n10271, n10272, 
        n10273, n10274, n10275, n10276, n10277, n10278, n10279, 
        n10280, n10281, n10282, n10283, n10284, n10285, n10286, 
        n10287, n10288, n10289, n10290, n10291, n10292, n10293, 
        n10294, n10295, n10296, n10297, n10298, n10299, n10300, 
        n10301, n10302, n10303, n10304, n10305, n10306, n10307, 
        n10308, n10309, n10310, n10311, n10312, n10313, n10314, 
        n10315, n10316, n10317, n10318, n10319, n10320, n10321, 
        n10322, n10323, n10324, n10325, n10326, n10327, n10328, 
        n10329, n10330, n10331, n10332, n10333, n10334, n10335, 
        n10336, n10337, n10338, n10339, n10340, n10341, n10342, 
        n10343, n10344, n10345, n10346, n10347, n10348, n10349, 
        n10350, n10351, n10352, n10353, n10354, n10355, n10356, 
        n10357, n10358, n10359, n10360, n10361, n10362, n10363, 
        n10364, n10365, n10366, n10367, n10368, n10369, n10370, 
        n10371, n10372, n10373, n10374, n10375, n10376, n10377, 
        n10378, n10379, n10380, n10381, n10382, n10383, n10384, 
        n10385, n10386, n10387, n10388, n10389, n10390, n10391, 
        n10392, n10393, n10394, n10395, n10396, n10397, n10398, 
        n10399, n10400, n10401, n10402, n10403, n10404, n10405, 
        n10406, n10407, n10408, n10409, n10410, n10411, n10412, 
        n10413, n10414, n10415, n10416, n10417, n10418, n10419, 
        n10420, n10421, n10422, n10423, n10424, n10425, n10426, 
        n10427, n10428, n10429, n10430, n10431, n10432, n10433, 
        n10434, n10435, n10436, n10437, n10438, n10439, n10440, 
        n10441, n10442, n10443, n10444, n10445, n10446, n10447, 
        n10448, n10449, n10450, n10451, n10452, n10453, n10454, 
        n10455, n10488, n10489, n10490, n10835, n10836, n10837, 
        n10838, n10852, n10853, n10854, n10855, n10856, n10857, 
        n10858, n10859, n10860, n10861, n10862, n10863, n10864, 
        n10865, n10866, n10867, n10868, n10869, n10870, n10871, 
        n10872, n10873, n10874, n10875, n10876, n10877, n10878, 
        n10879, n10880, n10881, n10882, n10883, n10884, n10885, 
        n10886, n10887, n10888, n10889, n10890, n10891, n10892, 
        n10893, n10894, n10895, n10896, n10897, n10898, n10899, 
        n10900, n10901, n10902, n10903, n10904, n10905, n10906, 
        n10907, n10908, n10909, n10910, n10911, n10912, n10913, 
        n10914, n10915, n10916, n10917, n10918, n10919, n10920, 
        n10921, n10922, n10923, n10924, n10925, n10926, n10927, 
        n10928, n10929, n10930, n10931, n10932, n10933, n10934, 
        n10935, n10936, n10937, n10938, n10939, n10940, n10941, 
        n10942, n10943, n10944, n10945, n10946, n10947, n10948, 
        n10949, n10950, n10951, n10952, n10953, n10954, n10955, 
        n10956, n10957, n10958, n10959, n10960, n10961, n10962, 
        n10963, n10964, n10965, n10966, n10967, n10968, n10969, 
        n10970, n10971, n10972, n10973, n10974, n10975, n10976, 
        n10977, n10978, n10979, n10980, n10981, n10982, n10983, 
        n10984, n10985, n10986, n10987, n10988, n10989, n10990, 
        n10991, n10992, n10993, n10994, n10995, n10996, n10997, 
        n10998, n10999, n11000, n11001, n11002, n11003, n11004, 
        n11005, n11006, n11007, n11008, n11009, n11010, n11011, 
        n11012, n11013, n11014, n11015, n11016, n11017, n11018, 
        n11019, n11020, n11021, n11022, n11023, n11024, n11025, 
        n11026, n11027, n11028, n11029, n11030, n11031, n11032, 
        n11033, n11034, n11035, n11036, n11037, n11038, n11039, 
        n11040, n11041, n11042, n11043, n11044, n11045, n11046, 
        n11047, n11048, n11049, n11050, n11051, n11052, n11053, 
        n11054, n11055, n11056, n11057, n11058, n11059, n11060, 
        n11061, n11062, n11063, n11064, n11065, n11066, n11067, 
        n11068, n11069, n11070, n11071, n11072, n11073, n11074, 
        n11075, n11076, n11077, n11078, n11079, n11080, n11081, 
        n11082, n11083, n11084, n11085, n11086, n11087, n11088, 
        n11089, n11090, n11091, n11092, n11093, n11094, n11095, 
        n11096, n11097, n11098, n11099, n11100, n11101, n11102, 
        n11103, n11104, n11105, n11106, n11107, n11108, n11109, 
        n11110, n11111, n11112, n11113, n11114, n11115, n11116, 
        n11117, n11118, n11119, n11120, n11121, n11122, n11123, 
        n11124, n11125, n11126, n11127, n11128, n11129, n11130, 
        n11131, n11132, n11133, n11134, n11135, n11136, n11137, 
        n11138, n11139, n11140, n11141, n11142, n11143, n11144, 
        n11145, n11146, n11147, n11148, n11149, n11150, n11151, 
        n11152, n11153, n11154, n11155, n11156, n11157, n11158, 
        n11159, n11160, n11161, n11162, n11163, n11164, n11165, 
        n11166, n11167, n11168, n11169, n11170, n11171, n11172, 
        n11173, n11174, n11175, n11176, n11177, n11178, n11179, 
        n11180, n11181, n11182, n11183, n11184, n11185, n11186, 
        n11187, n11188, n11189, n11190, n11191, n11192, n11193, 
        n11194, n11195, n11196, n11197, n11198, n11199, n11200, 
        n11201, n11202, n11203, n11204, n11205, n11206, n11207, 
        n11208, n11209, n11210, n11211, n11212, n11213, n11214, 
        n11215, n11216, n11217, n11218, n11219, n11220, n11221, 
        n11222, n11223, n11224, n11225, n11226, n11227, n11228, 
        n11229, n11230, n11231, n11232, n11233, n11234, n11235, 
        n11236, n11237, n11238, n11239, n11240, n11241, n11242, 
        n11243, n11244, n11245, n11246, n11247, n11248, n11249, 
        n11250, n11251, n11252, n11253, n11254, n11255, n11256, 
        n11257, n11258, n11259, n11260, n11261, n11262, n11263, 
        n11264, n11265, n11266, n11267, n11268, n11269, n11270, 
        n11271, n11272, n11273, n11274, n11275, n11276, n11277, 
        n11278, n11279, n11280, n11281, n11282, n11283, n11284, 
        n11285, n11286, n11287, n11288, n11289, n11290, n11291, 
        n11292, n11293, n11294, n11295, n11296, n11297, n11298, 
        n11299, n11300, n11301, n11302, n11303, n11304, n11305, 
        n11306, n11307, n11308, n11309, n11310, n11311, n11312, 
        n11313, n11314, n11315, n11316, n11317, n11318, n11319, 
        n11320, n11321, n11322, n11323, n11324, n11325, n11326, 
        n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
        n11334, n11335, n11336, n11337, n11338, n11339, n11340, 
        n11341, n11342, n11343, n11344, n11345, n11346, n11347, 
        n11348, n11349, n11350, n11351, n11352, n11353, n11354, 
        n11355, n11356, n11357, n11358, n11359, n11360, n11361, 
        n11362, n11363, n11364, n11365, n11366, n11367, n11368, 
        n11369, n11370, n11371, n11372, n11373, n11374, n11375, 
        n11376, n11377, n11378, n11379, n11380, n11381, n11382, 
        n11383, n11384, n11385, n11386, n11387, n11388, n11389, 
        n11390, n11391, n11392, n11393, n11394, n11395, n11396, 
        n11397, n11398, n11399, n11400, n11401, n11402, n11403, 
        n11404, n11405, n11406, n11407, n11408, n11409, n11410, 
        n11411, n11412, n11413, n11414, n11415, n11416, n11417, 
        n11418, n11419, n11420, n11421, n11422, n11423, n11424, 
        n11425, n11426, n11427, n11428, n11429, n11430, n11431, 
        n11432, n11433, n11434, n11435, n11436, n11437, n11438, 
        n11439, n11440, n11441, n11442, n11443, n11444, n11445, 
        n11446, n11447, n11448, n11449, n11450, n11451, n11452, 
        n11453, n11454, n11455, n11456, n11457, n11458, n11459, 
        n11460, n11461, n11462, n11463, n11464, n11465, n11466, 
        n11467, n11468, n11469, n11470, n11471, n11472, n11473, 
        n11474, n11475, n11476, n11477, n11478, n11479, n11480, 
        n11481, n11482, n11483, n11484, n11485, n11486, n11487, 
        n11488, n11489, n11490, n11491, n11492, n11493, n11494, 
        n11495, n11496, n11497, n11498, n11499, n11500, n11501, 
        n11502, n11503, n11504, n11505, n11506, n11507, n11508, 
        n11509, n11510, n11511, n11512, n11513, n11514, n11515, 
        n11516, n11517, n11518, n11519, n11520, n11521, n11522, 
        n11523, n11524, n11525, n11526, n11527, n11528, n11529, 
        n11530, n11531, n11532, n11533, n11534, n11535, n11536, 
        n11537, n11538, n11539, n11540, n11541, n11542, n11543, 
        n11544, n11545, n11546, n11547, n11548, n11549, n11550, 
        n11551, n11552, n11553, n11554, n11555, n11556, n11557, 
        n11558, n11559, n11560, n11561, n11562, n11563, n11564, 
        n11565, n11566, n11567, n11568, n11569, n11570, n11571, 
        n11572, n11573, n11574, n11575, n11576, n11577, n11578, 
        n11579, n11580, n11581, n11582, n11583, n11584, n11585, 
        n11586, n11587, n11588, n11589, n11590, n11591, n11592, 
        n11593, n11594, n11595, n11596, n11597, n11598, n11599, 
        n11600, n11601, n11602, n11603, n11604, n11605, n11606, 
        n11607, n11608, n11609, n11610, n11611, n11612, n11613, 
        n11614, n11615, n11616, n11617, n11618, n11619, n11620, 
        n11622, n11623, n11624, n11625, n11626, n11627, n11628, 
        n11629, n11630, n11631, n11632, n11633, n11634, n11635, 
        n11636, n11637, n11638, n11639, n11640, n11641, n11642, 
        n11643, n11644, n11645, n11646, n11647, n11648, n11649, 
        n11650, n11651, n11652, n11653, n11654, n11655, n11656, 
        n11657, n11658, n11659, n11660, n11661, n11662, n11663, 
        n11664, n11665, n11666, n11667, n11668, n11669, n11670, 
        n11671, n11672, n11673, n11674, n11675, n11676, n11677, 
        n11678, n11679, n11680, n11681, n11682, n11683, n11684, 
        n11685, n11686, n11687, n11688, n11689, n11690, n11691, 
        n11692, n11693, n11694, n11695, n11696, n11697, n11698, 
        n11699, n11700, n11701, n11702, n11703, n11704, n11705, 
        n11707, n11708, n11709, n11710, n11711, n11712, n11713, 
        n11714, n11715, n11716, n11717, n11718, n11719, n11720, 
        n11721, n11722, n11723, n11724, n11725, n11726, n11727, 
        n11728, n11729, n11730, n11731, n11732, n11733, n11734, 
        n11735, n11736, n11737, n11738, n11739, n11740, n11741, 
        n11742, n11743, n11744, n11745, n11746, n11747, n11748, 
        n11749, n11750, n11751, n11752, n11753, n11754, n11755, 
        n11756, n11757, n11758, n11759, n11760, n11761, n11762, 
        n11763, n11764, n11765, n11766, n11767, n11768, n11769, 
        n11770, n11771, n11772, n11773, n11774, n11775, n11776, 
        n11777, n11778, n11779, n11780, n11781, n11782, n11783, 
        n11784, n11785, n11786, n11787, n11788, n11789, n11790, 
        n11791, n11792, n11793, n11794, n11795, n11796, n11797, 
        n11798, n11799, n11800, n11801, n11802, n11803, n11804, 
        n11805, n11806, n11807, n11808, n11809, n11810, n11811, 
        n11812, n11813, n11814, n11815, n11816, n11817, n11818, 
        n11819, n11820, n11821, n11822, n11823, n11824, n11825, 
        n11826, n11827, n11828, n11829, n11830, n11831, n11832, 
        n11833, n11834, n11835, n11836, n11837, n11838, n11839, 
        n11840, n11841, n11842, n11843, n11844, n11845, n11846, 
        n11847, n11848, n11849, n11850, n11851, n11852, n11853, 
        n11854, n11855, n11856, n11857, n11858, n11859, n11860, 
        n11861, n11862, n11863, n11864, n11865, n12080, n12081, 
        n12082, n12083, n12084, n12085, n12086, n12087, n12088, 
        n12089, n12090, n12091, n12092, n12093, n12094, n12095, 
        n12096, n12097, n12098, n12099, n12100, n12101, n12102, 
        n12103, n12104, n12105, n12106, n12107, n12108, n12109, 
        n12110, n12111, n12112, n12113, n12114, n12115, n12116, 
        n12117, n12118, n12120, n12121, n12122, n12123, n12124, 
        n12125, n12126, n12127, n12128, n12129, n12130, n12131, 
        n12132, n12133, n12134, n12135, n12136, n12137, n12138, 
        n12139, n12140;
    
    assign mipi_resetn_o = hdmi_resetn_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_resetn_o = PllLocked[1] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign DdrCtrl_AID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[31] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[30] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[29] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[28] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[27] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[26] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[25] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[24] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[3] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[2] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[1] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[2] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ABURST_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ABURST_0[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[15] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[14] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[13] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[12] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[11] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[10] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[9] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[8] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[7] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[6] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[5] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[4] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[3] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[2] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[1] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_BREADY_0 = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lcd_pwm = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[4] = hdmi_txc_o[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[3] = hdmi_txc_o[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[2] = hdmi_txc_o[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[1] = hdmi_txc_o[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi0_scl_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi0_scl_oe = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi0_sda_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi0_sda_oe = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi1_scl_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi1_scl_oe = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi1_sda_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi1_sda_oe = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_trig_o[1] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_trig_o[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_RSTN_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_DPHY_RSTN_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_VC_ENA_o[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_VC_ENA_o[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_VC_ENA_o[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_VC_ENA_o[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_LANES_o[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_0_LANES_o[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_RSTN_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_DPHY_RSTN_o = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_VC_ENA_o[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_VC_ENA_o[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_VC_ENA_o[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_VC_ENA_o[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_LANES_o[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_LANES_o[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_rx_1_CLEAR = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_RREADY_0 = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign mipi_rx_0_CLEAR = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 LUT__13701 (.I0(\DdrCtrl_ARADDR_0[23] ), .I1(\DdrCtrl_AWADDR_0[23] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13701.LUTMASK = 16'hcaca;
    EFX_FF \Axi0ResetReg[2]~FF  (.D(\Axi0ResetReg[1] ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(270)
    defparam \Axi0ResetReg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[1]~FF  (.D(\Axi0ResetReg[0] ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(270)
    defparam \Axi0ResetReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ResetShiftReg[0]~FF  (.D(\reduce_nand_9/n7 ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(231)
    defparam \ResetShiftReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[0]~FF  (.D(DdrInitDone), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(270)
    defparam \Axi0ResetReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_vsync~FF  (.D(w_XYCrop0_frame_vsync), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(r_XYCrop0_frame_vsync)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_vsync~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_vsync~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_vsync~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_vsync~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_vsync~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_vsync~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_vsync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[0]~FF  (.D(\w_XYCrop0_frame_Gray[0] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[0]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[0]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[0]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[0]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[0]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[0]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_href~FF  (.D(w_XYCrop0_frame_href), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(r_XYCrop0_frame_href)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_href~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_href~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_href~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_href~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_href~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_href~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_href~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_de~FF  (.D(w_XYCrop0_frame_de), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(r_XYCrop0_frame_de)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_de~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_de~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_de~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_de~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_de~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_de~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_de~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_rst_n~FF  (.D(\Axi0ResetReg[2] ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(r_hdmi_rst_n)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(532)
    defparam \r_hdmi_rst_n~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_rst_n~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_RSTN~FF  (.D(\ResetShiftReg[1] ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(DdrCtrl_RSTN)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(231)
    defparam \DdrCtrl_RSTN~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_RSTN~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_RSTN~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_RSTN~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_RSTN~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_RSTN~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_RSTN~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ResetShiftReg[1]~FF  (.D(\ResetShiftReg[0] ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(231)
    defparam \ResetShiftReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrInitDone~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n58 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(DdrInitDone)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \DdrInitDone~FF .CLK_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .CE_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .SR_POLARITY = 1'b0;
    defparam \DdrInitDone~FF .D_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .SR_SYNC = 1'b0;
    defparam \DdrInitDone~FF .SR_VALUE = 1'b0;
    defparam \DdrInitDone~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rc_hdmi_tx~FF  (.D(rc_hdmi_tx), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(rc_hdmi_tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \rc_hdmi_tx~FF .CLK_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .CE_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .SR_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .D_POLARITY = 1'b0;
    defparam \rc_hdmi_tx~FF .SR_SYNC = 1'b1;
    defparam \rc_hdmi_tx~FF .SR_VALUE = 1'b0;
    defparam \rc_hdmi_tx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[0]~FF  (.D(n927_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx0_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[0]~FF  (.D(n938_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx1_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[0]~FF  (.D(n949_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx2_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[0]~FF  (.D(n33_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_CFG_SEQ_START~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n89 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(DdrCtrl_CFG_SEQ_START)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(187)
    defparam \DdrCtrl_CFG_SEQ_START~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(187)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(151)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(151)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n57 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(187)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n56 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n55 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n54 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n53 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n52 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n51 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n50 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n49 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n48 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n47 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n46 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n45 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n44 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n43 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n42 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n41 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n40 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n39 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n38 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(DdrCtrl_RSTN), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(172)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16bit/n158 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/current_state[0]~FF  (.D(\u_i2c_timing_ctrl_16bit/n189 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/current_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(146)
    defparam \u_i2c_timing_ctrl_16bit/current_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF  (.D(\u_i2c_timing_ctrl_16bit/n159 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_ctrl_clk )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_ctrl_clk~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF  (.D(\u_i2c_timing_ctrl_16bit/n160 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_transfer_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_transfer_en~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[0]~FF  (.D(\u_i2c_timing_ctrl_16bit/n241 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[0]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[0]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16bit/n374 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF  (.D(\u_i2c_timing_ctrl_16bit/n383 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF  (.D(\u_i2c_timing_ctrl_16bit/n63 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16bit/n64 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cmos_sdat_OUT~FF  (.D(\u_i2c_timing_ctrl_16bit/n369 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(cmos_sdat_OUT)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \cmos_sdat_OUT~FF .CLK_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .CE_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_POLARITY = 1'b0;
    defparam \cmos_sdat_OUT~FF .D_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_SYNC = 1'b0;
    defparam \cmos_sdat_OUT~FF .SR_VALUE = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF  (.D(\u_i2c_timing_ctrl_16bit/n157 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF  (.D(\u_i2c_timing_ctrl_16bit/n156 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF  (.D(\u_i2c_timing_ctrl_16bit/n155 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF  (.D(\u_i2c_timing_ctrl_16bit/n154 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF  (.D(\u_i2c_timing_ctrl_16bit/n153 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF  (.D(\u_i2c_timing_ctrl_16bit/n152 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF  (.D(\u_i2c_timing_ctrl_16bit/n151 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF  (.D(\u_i2c_timing_ctrl_16bit/n150 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF  (.D(\u_i2c_timing_ctrl_16bit/n149 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF  (.D(\u_i2c_timing_ctrl_16bit/n148 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF  (.D(\u_i2c_timing_ctrl_16bit/n147 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF  (.D(\u_i2c_timing_ctrl_16bit/n146 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF  (.D(\u_i2c_timing_ctrl_16bit/n145 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF  (.D(\u_i2c_timing_ctrl_16bit/n144 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF  (.D(\u_i2c_timing_ctrl_16bit/n143 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/clk_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(119)
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/clk_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/current_state[1]~FF  (.D(\u_i2c_timing_ctrl_16bit/n188 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/current_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(146)
    defparam \u_i2c_timing_ctrl_16bit/current_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/current_state[2]~FF  (.D(\u_i2c_timing_ctrl_16bit/n187 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/current_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(146)
    defparam \u_i2c_timing_ctrl_16bit/current_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/current_state[3]~FF  (.D(\u_i2c_timing_ctrl_16bit/n186 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/current_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(146)
    defparam \u_i2c_timing_ctrl_16bit/current_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/current_state[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/current_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[1]~FF  (.D(\u_i2c_timing_ctrl_16bit/n240 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[1]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[1]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[2]~FF  (.D(\u_i2c_timing_ctrl_16bit/n239 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[2]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[2]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[3]~FF  (.D(\u_i2c_timing_ctrl_16bit/n238 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[3]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[3]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[4]~FF  (.D(\u_i2c_timing_ctrl_16bit/n237 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[4]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[4]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[5]~FF  (.D(\u_i2c_timing_ctrl_16bit/n236 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[5]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[5]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[6]~FF  (.D(\u_i2c_timing_ctrl_16bit/n235 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[6]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[6]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[7]~FF  (.D(\u_i2c_timing_ctrl_16bit/n234 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[7]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[7]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[8]~FF  (.D(\u_i2c_timing_ctrl_16bit/n233 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(173)
    defparam \i2c_config_index[8]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[8]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[8]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[8]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[8]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[8]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF  (.D(\u_i2c_timing_ctrl_16bit/n373 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF  (.D(\u_i2c_timing_ctrl_16bit/n372 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF  (.D(\u_i2c_timing_ctrl_16bit/n371 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF  (.D(\u_i2c_timing_ctrl_16bit/n382 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF  (.D(\u_i2c_timing_ctrl_16bit/n381 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF  (.D(\u_i2c_timing_ctrl_16bit/n380 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF  (.D(\u_i2c_timing_ctrl_16bit/n379 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF  (.D(\u_i2c_timing_ctrl_16bit/n378 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF  (.D(\u_i2c_timing_ctrl_16bit/n377 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF  (.D(\u_i2c_timing_ctrl_16bit/n376 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/i2c_wdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(322)
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/i2c_wdata[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF  (.D(\u_i2c_timing_ctrl_16bit/n62 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF  (.D(\u_i2c_timing_ctrl_16bit/n61 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF  (.D(\u_i2c_timing_ctrl_16bit/n60 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF  (.D(\u_i2c_timing_ctrl_16bit/n59 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF  (.D(\u_i2c_timing_ctrl_16bit/n58 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF  (.D(\u_i2c_timing_ctrl_16bit/n57 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF  (.D(\u_i2c_timing_ctrl_16bit/n56 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF  (.D(\u_i2c_timing_ctrl_16bit/n55 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF  (.D(\u_i2c_timing_ctrl_16bit/n54 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF  (.D(\u_i2c_timing_ctrl_16bit/n53 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF  (.D(\u_i2c_timing_ctrl_16bit/n52 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF  (.D(\u_i2c_timing_ctrl_16bit/n51 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF  (.D(\u_i2c_timing_ctrl_16bit/n50 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF  (.D(\u_i2c_timing_ctrl_16bit/n49 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF  (.D(\u_i2c_timing_ctrl_16bit/n48 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF  (.D(\u_i2c_timing_ctrl_16bit/n47 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF  (.D(\u_i2c_timing_ctrl_16bit/n46 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF  (.D(\u_i2c_timing_ctrl_16bit/n45 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF  (.D(\u_i2c_timing_ctrl_16bit/n44 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF  (.D(\u_i2c_timing_ctrl_16bit/n43 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF  (.D(\u_i2c_timing_ctrl_16bit/n42 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF  (.D(\u_i2c_timing_ctrl_16bit/n41 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF  (.D(\u_i2c_timing_ctrl_16bit/n40 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF  (.D(\u_i2c_timing_ctrl_16bit/n39 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF  (.D(\u_i2c_timing_ctrl_16bit/n38 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16bit/delay_cnt[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(69)
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16bit/delay_cnt[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF  (.D(\u_Sensor_Image_XYCrop_0/n42 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF  (.D(\u_Sensor_Image_XYCrop_0/n43 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF  (.D(\u_Sensor_Image_XYCrop_0/n44 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_in_href_r~FF  (.D(cmos_href), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_Sensor_Image_XYCrop_0/image_in_href_r )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \u_Sensor_Image_XYCrop_0/image_in_href_r~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_in_href_r~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_in_href_r~FF .SR_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_in_href_r~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_in_href_r~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_in_href_r~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_in_href_r~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF  (.D(\u_Sensor_Image_XYCrop_0/n53 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_de~FF  (.D(1'b1), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(w_XYCrop0_frame_de)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_de~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_de~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_de~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_de~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_de~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_de~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_de~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF  (.D(\u_Sensor_Image_XYCrop_0/n45 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF  (.D(\u_Sensor_Image_XYCrop_0/n46 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[5]~FF  (.D(cmos_data[5]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[5]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[5]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[5]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[5]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[5]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[5]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF  (.D(\u_Sensor_Image_XYCrop_0/n47 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF  (.D(\u_Sensor_Image_XYCrop_0/n48 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF  (.D(\u_Sensor_Image_XYCrop_0/image_xpos[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF .D_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[3]~FF  (.D(cmos_data[3]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[3]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[3]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[3]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[3]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[3]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[3]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF  (.D(\u_Sensor_Image_XYCrop_0/n49 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF  (.D(\u_Sensor_Image_XYCrop_0/n50 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[4]~FF  (.D(cmos_data[4]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[4]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[4]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[4]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[4]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF  (.D(\u_Sensor_Image_XYCrop_0/n51 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_href~FF  (.D(\u_Sensor_Image_XYCrop_0/w_image_out_href ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(w_XYCrop0_frame_href)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(127)
    defparam \w_XYCrop0_frame_href~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_href~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_href~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_href~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_href~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_href~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_href~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF  (.D(\u_Sensor_Image_XYCrop_0/n52 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(cmos_vsync), .Q(\u_Sensor_Image_XYCrop_0/image_ypos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(99)
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_ypos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[6]~FF  (.D(cmos_data[6]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[6]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[6]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[6]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[6]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[6]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[6]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[7]~FF  (.D(cmos_data[7]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[7]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[7]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[7]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[7]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[7]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[7]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[2]~FF  (.D(cmos_data[2]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[2]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[2]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[2]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[2]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[2]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[2]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[1]~FF  (.D(cmos_data[1]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[1]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[1]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[1]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[1]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[1]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[1]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_Gray[0]~FF  (.D(cmos_data[0]), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(\w_XYCrop0_frame_Gray[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_Gray[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[0]~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[0]~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_Gray[0]~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_Gray[0]~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_Gray[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_XYCrop0_frame_vsync~FF  (.D(cmos_vsync), .CE(1'b1), .CLK(\cmos_pclk~O ), 
           .SR(1'b0), .Q(w_XYCrop0_frame_vsync)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(79)
    defparam \w_XYCrop0_frame_vsync~FF .CLK_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_vsync~FF .CE_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_vsync~FF .SR_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_vsync~FF .D_POLARITY = 1'b1;
    defparam \w_XYCrop0_frame_vsync~FF .SR_SYNC = 1'b1;
    defparam \w_XYCrop0_frame_vsync~FF .SR_VALUE = 1'b0;
    defparam \w_XYCrop0_frame_vsync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF  (.D(n463), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF  (.D(n4419), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF  (.D(n4417), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF  (.D(n4415), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF  (.D(n4413), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF  (.D(n4411), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF  (.D(n4409), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF  (.D(n4407), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF  (.D(n4405), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF  (.D(n4403), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF  (.D(n4402), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(cmos_href), .Q(\u_Sensor_Image_XYCrop_0/image_xpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(115)
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF .D_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF .SR_SYNC = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF .SR_VALUE = 1'b0;
    defparam \u_Sensor_Image_XYCrop_0/image_xpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[1]~FF  (.D(\w_XYCrop0_frame_Gray[1] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[1]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[1]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[1]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[1]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[1]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[1]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[2]~FF  (.D(\w_XYCrop0_frame_Gray[2] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[2]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[2]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[2]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[2]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[2]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[2]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[3]~FF  (.D(\w_XYCrop0_frame_Gray[3] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[3]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[3]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[3]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[3]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[3]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[3]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[4]~FF  (.D(\w_XYCrop0_frame_Gray[4] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[4]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[4]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[4]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[4]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[4]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[4]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[5]~FF  (.D(\w_XYCrop0_frame_Gray[5] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[5]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[5]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[5]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[5]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[6]~FF  (.D(\w_XYCrop0_frame_Gray[6] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[6]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[6]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[6]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[6]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_XYCrop0_frame_Gray[7]~FF  (.D(\w_XYCrop0_frame_Gray[7] ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\r_XYCrop0_frame_Gray[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(384)
    defparam \r_XYCrop0_frame_Gray[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[7]~FF .SR_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[7]~FF .D_POLARITY = 1'b1;
    defparam \r_XYCrop0_frame_Gray[7]~FF .SR_SYNC = 1'b1;
    defparam \r_XYCrop0_frame_Gray[7]~FF .SR_VALUE = 1'b0;
    defparam \r_XYCrop0_frame_Gray[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \axi4_awar_mux/rs_req[0]~FF  (.D(\axi4_awar_mux/n50 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\axi4_awar_mux/rs_req[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\AXI4_AWARMux.v(105)
    defparam \axi4_awar_mux/rs_req[0]~FF .CLK_POLARITY = 1'b1;
    defparam \axi4_awar_mux/rs_req[0]~FF .CE_POLARITY = 1'b1;
    defparam \axi4_awar_mux/rs_req[0]~FF .SR_POLARITY = 1'b0;
    defparam \axi4_awar_mux/rs_req[0]~FF .D_POLARITY = 1'b1;
    defparam \axi4_awar_mux/rs_req[0]~FF .SR_SYNC = 1'b1;
    defparam \axi4_awar_mux/rs_req[0]~FF .SR_VALUE = 1'b0;
    defparam \axi4_awar_mux/rs_req[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWREADY_0~FF  (.D(DdrCtrl_ATYPE_0), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(\axi4_awar_mux/n131 ), .Q(DdrCtrl_AWREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\AXI4_AWARMux.v(105)
    defparam \DdrCtrl_AWREADY_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWREADY_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWREADY_0~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWREADY_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWREADY_0~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AWREADY_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWREADY_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AVALID_0~FF  (.D(\axi4_awar_mux/n52 ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\AXI4_AWARMux.v(105)
    defparam \DdrCtrl_AVALID_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AVALID_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AVALID_0~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AVALID_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AVALID_0~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AVALID_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AVALID_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ATYPE_0~FF  (.D(\axi4_awar_mux/n55 ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_ATYPE_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\AXI4_AWARMux.v(105)
    defparam \DdrCtrl_ATYPE_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_ATYPE_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARREADY_0~FF  (.D(DdrCtrl_ATYPE_0), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(\axi4_awar_mux/n131 ), .Q(DdrCtrl_ARREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\AXI4_AWARMux.v(105)
    defparam \DdrCtrl_ARREADY_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARREADY_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARREADY_0~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_ARREADY_0~FF .D_POLARITY = 1'b0;
    defparam \DdrCtrl_ARREADY_0~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ARREADY_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARREADY_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \axi4_awar_mux/rs_req[1]~FF  (.D(\axi4_awar_mux/n49 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\axi4_awar_mux/rs_req[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\AXI4_AWARMux.v(105)
    defparam \axi4_awar_mux/rs_req[1]~FF .CLK_POLARITY = 1'b1;
    defparam \axi4_awar_mux/rs_req[1]~FF .CE_POLARITY = 1'b1;
    defparam \axi4_awar_mux/rs_req[1]~FF .SR_POLARITY = 1'b0;
    defparam \axi4_awar_mux/rs_req[1]~FF .D_POLARITY = 1'b1;
    defparam \axi4_awar_mux/rs_req[1]~FF .SR_SYNC = 1'b1;
    defparam \axi4_awar_mux/rs_req[1]~FF .SR_VALUE = 1'b0;
    defparam \axi4_awar_mux/rs_req[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wframe_index_last[1]~FF  (.D(\u_axi4_ctrl_0/n119 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_wframe_index_last[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(154)
    defparam \u_axi4_ctrl_0/r_wframe_index_last[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[23]~FF  (.D(\u_axi4_ctrl_0/n116 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_ARADDR_0[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(154)
    defparam \DdrCtrl_ARADDR_0[23]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[23]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[23]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_ARADDR_0[23]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[23]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ARADDR_0[23]~FF .SR_VALUE = 1'b1;
    defparam \DdrCtrl_ARADDR_0[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[22]~FF  (.D(\u_axi4_ctrl_0/n117 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_ARADDR_0[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(154)
    defparam \DdrCtrl_ARADDR_0[22]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[22]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[22]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_ARADDR_0[22]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[22]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ARADDR_0[22]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wframe_index_last[0]~FF  (.D(\u_axi4_ctrl_0/n120 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_wframe_index_last[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(154)
    defparam \u_axi4_ctrl_0/r_wframe_index_last[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_index_last[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rs_w[0]~FF  (.D(\u_axi4_ctrl_0/n265 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/rs_w[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rs_w[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rs_w[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rs_w[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rs_w[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rs_w[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rs_w[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rs_w[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[0]~FF  (.D(\u_axi4_ctrl_0/n290 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[0]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[0]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[0]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[0]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[0]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wframe_sync[0]~FF  (.D(r_XYCrop0_frame_vsync), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_wframe_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/r_wframe_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_sync[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_sync[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_w_eof[0]~FF  (.D(\u_axi4_ctrl_0/n291 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/rc_w_eof[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_w_eof[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_w_eof[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_w_eof[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rc_w_eof[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_w_eof[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rc_w_eof[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_w_eof[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWVALID_0~FF  (.D(\u_axi4_ctrl_0/n258 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AWVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWVALID_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWVALID_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWVALID_0~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWVALID_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWVALID_0~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWVALID_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWVALID_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_WVALID_0~FF  (.D(\u_axi4_ctrl_0/n260 ), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_WVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_WVALID_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_WVALID_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_WVALID_0~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_WVALID_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_WVALID_0~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_WVALID_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_WVALID_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[0]~FF  (.D(\u_axi4_ctrl_0/n346 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_weof_pending~FF  (.D(\u_axi4_ctrl_0/n267 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_weof_pending )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/r_weof_pending~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_weof_pending~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_weof_pending~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_weof_pending~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_weof_pending~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/r_weof_pending~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_weof_pending~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wframe_inc~FF  (.D(\u_axi4_ctrl_0/n266 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_wframe_inc )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/r_wframe_inc~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_inc~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_inc~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_inc~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_inc~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_inc~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_inc~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_wfifo_we[0]~FF  (.D(\u_axi4_ctrl_0/n2649 ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), .Q(\u_axi4_ctrl_0/rc_wfifo_we[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/rc_wfifo_we[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rframe_vsync_dly~FF  (.D(lcd_vs), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/rframe_vsync_dly )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(340)
    defparam \u_axi4_ctrl_0/rframe_vsync_dly~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rframe_vsync_dly~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rframe_vsync_dly~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rframe_vsync_dly~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rframe_vsync_dly~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rframe_vsync_dly~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rframe_vsync_dly~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_cnt[1]~FF  (.D(\u_axi4_ctrl_0/n1074 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/n2551 ), .Q(\u_axi4_ctrl_0/rfifo_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(360)
    defparam \u_axi4_ctrl_0/rfifo_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_cnt[0]~FF  (.D(\u_axi4_ctrl_0/n1075 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/n2551 ), .Q(\u_axi4_ctrl_0/rfifo_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(360)
    defparam \u_axi4_ctrl_0/rfifo_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_rst~FF  (.D(\u_axi4_ctrl_0/equal_138/n9 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_axi4_ctrl_0/rfifo_rst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(375)
    defparam \u_axi4_ctrl_0/rfifo_rst~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_rst~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_rst~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_rst~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_rst~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_rst~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_rst~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rfifo_rst~FF  (.D(\u_axi4_ctrl_0/w_rfifo_rst ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rfifo_rst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(411)
    defparam \u_axi4_ctrl_0/r_rfifo_rst~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rfifo_rst~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF  (.D(\u_axi4_ctrl_0/n2670 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst_rclk ), 
           .Q(\u_axi4_ctrl_0/rc_rfifo_rd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(427)
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF  (.D(\u_axi4_ctrl_0/w_rfifo_rst ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rfifo_rst_rclk )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(416)
    defparam \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rfifo_rst_rclk~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF  (.D(1'b1), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_inc~FF  (.D(\u_axi4_ctrl_0/equal_160/n3 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_rframe_inc )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(480)
    defparam \u_axi4_ctrl_0/r_rframe_inc~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_inc~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_inc~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_inc~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_inc~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_inc~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_inc~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF  (.D(\u_axi4_ctrl_0/n1730 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rd_state.S_READ_IDLE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(553)
    defparam \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_IDLE~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF  (.D(\u_axi4_ctrl_0/select_190/Select_1/n3 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rd_state.S_READ_ADDR )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(553)
    defparam \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_ADDR~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF  (.D(\u_axi4_ctrl_0/n1732 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rd_state.S_READ_DATA )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(553)
    defparam \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rd_state.S_READ_DATA~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARVALID_0~FF  (.D(\u_axi4_ctrl_0/n1733 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(DdrCtrl_ARVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(553)
    defparam \DdrCtrl_ARVALID_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARVALID_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARVALID_0~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARVALID_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARVALID_0~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARVALID_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARVALID_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rd_pend~FF  (.D(\u_axi4_ctrl_0/n1734 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\u_axi4_ctrl_0/r_rd_pend )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(553)
    defparam \u_axi4_ctrl_0/r_rd_pend~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rd_pend~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rd_pend~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rd_pend~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rd_pend~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/r_rd_pend~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rd_pend~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wenb~FF  (.D(DdrCtrl_RVALID_0), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/rfifo_wenb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(605)
    defparam \u_axi4_ctrl_0/rfifo_wenb~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wenb~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wenb~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wenb~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wenb~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wenb~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wenb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[3]~FF  (.D(DdrCtrl_RDATA_0[3]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[2]~FF  (.D(DdrCtrl_RDATA_0[2]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[1]~FF  (.D(DdrCtrl_RDATA_0[1]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[0]~FF  (.D(DdrCtrl_RDATA_0[0]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rs_w[1]~FF  (.D(\u_axi4_ctrl_0/n264 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/rs_w[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rs_w[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rs_w[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rs_w[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rs_w[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rs_w[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rs_w[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rs_w[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[22]~FF  (.D(\u_axi4_ctrl_0/n2777 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(154)
    defparam \DdrCtrl_AWADDR_0[22]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[22]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[22]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[22]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[22]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AWADDR_0[22]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_w_rst~FF  (.D(\u_axi4_ctrl_0/n256 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_w_rst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/r_w_rst~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_w_rst~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_w_rst~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_w_rst~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_w_rst~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/r_w_rst~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_w_rst~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[1]~FF  (.D(\u_axi4_ctrl_0/n289 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[1]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[1]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[1]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[1]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[1]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[2]~FF  (.D(\u_axi4_ctrl_0/n288 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[2]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[2]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[2]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[2]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[2]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[3]~FF  (.D(\u_axi4_ctrl_0/n287 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[3]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[3]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[3]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[3]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[3]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[4]~FF  (.D(\u_axi4_ctrl_0/n286 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[4]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[4]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[4]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[4]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[4]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[5]~FF  (.D(\u_axi4_ctrl_0/n285 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[5]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[5]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[5]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[5]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[5]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[6]~FF  (.D(\u_axi4_ctrl_0/n284 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[6]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[6]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[6]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[6]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[6]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[7]~FF  (.D(\u_axi4_ctrl_0/n283 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[7]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[7]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[7]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[7]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[7]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[8]~FF  (.D(\u_axi4_ctrl_0/n282 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[8]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[8]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[8]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[8]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[8]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[9]~FF  (.D(\u_axi4_ctrl_0/n281 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[9]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[9]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[9]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[9]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[9]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[10]~FF  (.D(\u_axi4_ctrl_0/n280 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[10]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[10]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[10]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[10]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[10]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[11]~FF  (.D(\u_axi4_ctrl_0/n279 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[11]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[11]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[11]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[11]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[11]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[12]~FF  (.D(\u_axi4_ctrl_0/n278 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[12]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[12]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[12]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[12]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[12]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[13]~FF  (.D(\u_axi4_ctrl_0/n277 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[13]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[13]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[13]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[13]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[13]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[14]~FF  (.D(\u_axi4_ctrl_0/n276 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[14]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[14]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[14]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[14]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[14]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[15]~FF  (.D(\u_axi4_ctrl_0/n275 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[15]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[15]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[15]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[15]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[15]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[16]~FF  (.D(\u_axi4_ctrl_0/n274 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[16]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[16]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[16]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[16]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[16]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[17]~FF  (.D(\u_axi4_ctrl_0/n273 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[17]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[17]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[17]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[17]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[17]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[18]~FF  (.D(\u_axi4_ctrl_0/n272 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[18]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[18]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[18]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[18]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[18]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[19]~FF  (.D(\u_axi4_ctrl_0/n271 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[19]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[19]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[19]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[19]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[19]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[20]~FF  (.D(\u_axi4_ctrl_0/n270 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[20]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[20]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[20]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[20]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[20]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[21]~FF  (.D(\u_axi4_ctrl_0/n269 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \DdrCtrl_AWADDR_0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[21]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[21]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[21]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[21]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_AWADDR_0[21]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wframe_sync[1]~FF  (.D(\u_axi4_ctrl_0/r_wframe_sync[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl_0/r_wframe_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/r_wframe_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_sync[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wframe_sync[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wframe_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[1]~FF  (.D(\u_axi4_ctrl_0/n345 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[2]~FF  (.D(\u_axi4_ctrl_0/n344 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[3]~FF  (.D(\u_axi4_ctrl_0/n343 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[4]~FF  (.D(\u_axi4_ctrl_0/n342 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[5]~FF  (.D(\u_axi4_ctrl_0/n341 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[6]~FF  (.D(\u_axi4_ctrl_0/n340 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_burst[7]~FF  (.D(\u_axi4_ctrl_0/n339 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rc_burst[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl_0/rc_burst[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_burst[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_burst[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF  (.D(\u_axi4_ctrl_0/n766 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF  (.D(\u_axi4_ctrl_0/n765 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF  (.D(\u_axi4_ctrl_0/n764 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF  (.D(\u_axi4_ctrl_0/n763 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF  (.D(\u_axi4_ctrl_0/n762 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF  (.D(\u_axi4_ctrl_0/n761 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF  (.D(\u_axi4_ctrl_0/n760 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF  (.D(\u_axi4_ctrl_0/n759 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF  (.D(\u_axi4_ctrl_0/n758 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF  (.D(\u_axi4_ctrl_0/n757 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF  (.D(\u_axi4_ctrl_0/n756 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF  (.D(\u_axi4_ctrl_0/n755 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF  (.D(\u_axi4_ctrl_0/n754 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF  (.D(\u_axi4_ctrl_0/n753 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF  (.D(\u_axi4_ctrl_0/n752 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF  (.D(\u_axi4_ctrl_0/n751 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF  (.D(\u_axi4_ctrl_0/n750 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF  (.D(\u_axi4_ctrl_0/n749 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF  (.D(\u_axi4_ctrl_0/n748 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF  (.D(\u_axi4_ctrl_0/n747 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF  (.D(\u_axi4_ctrl_0/n746 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF  (.D(\u_axi4_ctrl_0/n745 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF  (.D(\u_axi4_ctrl_0/n744 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF  (.D(\u_axi4_ctrl_0/n743 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF  (.D(\u_axi4_ctrl_0/n742 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF  (.D(\u_axi4_ctrl_0/n741 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF  (.D(\u_axi4_ctrl_0/n740 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF  (.D(\u_axi4_ctrl_0/n739 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF  (.D(\u_axi4_ctrl_0/n738 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF  (.D(\u_axi4_ctrl_0/n737 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF  (.D(\u_axi4_ctrl_0/n736 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF  (.D(\u_axi4_ctrl_0/n735 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF  (.D(\u_axi4_ctrl_0/n734 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF  (.D(\u_axi4_ctrl_0/n733 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF  (.D(\u_axi4_ctrl_0/n732 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF  (.D(\u_axi4_ctrl_0/n731 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF  (.D(\u_axi4_ctrl_0/n730 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF  (.D(\u_axi4_ctrl_0/n729 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF  (.D(\u_axi4_ctrl_0/n728 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF  (.D(\u_axi4_ctrl_0/n727 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF  (.D(\u_axi4_ctrl_0/n726 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF  (.D(\u_axi4_ctrl_0/n725 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF  (.D(\u_axi4_ctrl_0/n724 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF  (.D(\u_axi4_ctrl_0/n723 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF  (.D(\u_axi4_ctrl_0/n722 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF  (.D(\u_axi4_ctrl_0/n721 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF  (.D(\u_axi4_ctrl_0/n720 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF  (.D(\u_axi4_ctrl_0/n719 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF  (.D(\u_axi4_ctrl_0/n718 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF  (.D(\u_axi4_ctrl_0/n717 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF  (.D(\u_axi4_ctrl_0/n716 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF  (.D(\u_axi4_ctrl_0/n715 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF  (.D(\u_axi4_ctrl_0/n714 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF  (.D(\u_axi4_ctrl_0/n713 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF  (.D(\u_axi4_ctrl_0/n712 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF  (.D(\u_axi4_ctrl_0/n711 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF  (.D(\u_axi4_ctrl_0/n710 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF  (.D(\u_axi4_ctrl_0/n709 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF  (.D(\u_axi4_ctrl_0/n708 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF  (.D(\u_axi4_ctrl_0/n707 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF  (.D(\u_axi4_ctrl_0/n706 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF  (.D(\u_axi4_ctrl_0/n705 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF  (.D(\u_axi4_ctrl_0/n704 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF  (.D(\u_axi4_ctrl_0/n703 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF  (.D(\u_axi4_ctrl_0/n702 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF  (.D(\u_axi4_ctrl_0/n701 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF  (.D(\u_axi4_ctrl_0/n700 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF  (.D(\u_axi4_ctrl_0/n699 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF  (.D(\u_axi4_ctrl_0/n698 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF  (.D(\u_axi4_ctrl_0/n697 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF  (.D(\u_axi4_ctrl_0/n696 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF  (.D(\u_axi4_ctrl_0/n695 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF  (.D(\u_axi4_ctrl_0/n694 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF  (.D(\u_axi4_ctrl_0/n693 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF  (.D(\u_axi4_ctrl_0/n692 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF  (.D(\u_axi4_ctrl_0/n691 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF  (.D(\u_axi4_ctrl_0/n690 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF  (.D(\u_axi4_ctrl_0/n689 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF  (.D(\u_axi4_ctrl_0/n688 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF  (.D(\u_axi4_ctrl_0/n687 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF  (.D(\u_axi4_ctrl_0/n686 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF  (.D(\u_axi4_ctrl_0/n685 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF  (.D(\u_axi4_ctrl_0/n684 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF  (.D(\u_axi4_ctrl_0/n683 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF  (.D(\u_axi4_ctrl_0/n682 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF  (.D(\u_axi4_ctrl_0/n681 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF  (.D(\u_axi4_ctrl_0/n680 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF  (.D(\u_axi4_ctrl_0/n679 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF  (.D(\u_axi4_ctrl_0/n678 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF  (.D(\u_axi4_ctrl_0/n677 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF  (.D(\u_axi4_ctrl_0/n676 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF  (.D(\u_axi4_ctrl_0/n675 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF  (.D(\u_axi4_ctrl_0/n674 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF  (.D(\u_axi4_ctrl_0/n673 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF  (.D(\u_axi4_ctrl_0/n672 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF  (.D(\u_axi4_ctrl_0/n671 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF  (.D(\u_axi4_ctrl_0/n670 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF  (.D(\u_axi4_ctrl_0/n669 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF  (.D(\u_axi4_ctrl_0/n668 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF  (.D(\u_axi4_ctrl_0/n667 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF  (.D(\u_axi4_ctrl_0/n666 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF  (.D(\u_axi4_ctrl_0/n665 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF  (.D(\u_axi4_ctrl_0/n664 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF  (.D(\u_axi4_ctrl_0/n663 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF  (.D(\u_axi4_ctrl_0/n662 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF  (.D(\u_axi4_ctrl_0/n661 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF  (.D(\u_axi4_ctrl_0/n660 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF  (.D(\u_axi4_ctrl_0/n659 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF  (.D(\u_axi4_ctrl_0/n658 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF  (.D(\u_axi4_ctrl_0/n657 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF  (.D(\u_axi4_ctrl_0/n656 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF  (.D(\u_axi4_ctrl_0/n655 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF  (.D(\u_axi4_ctrl_0/n654 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF  (.D(\u_axi4_ctrl_0/n653 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF  (.D(\u_axi4_ctrl_0/n652 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF  (.D(\u_axi4_ctrl_0/n651 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF  (.D(\u_axi4_ctrl_0/n650 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF  (.D(\u_axi4_ctrl_0/n649 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF  (.D(\u_axi4_ctrl_0/n648 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF  (.D(\u_axi4_ctrl_0/n647 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_wfifo_wdata[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_wfifo_wdata[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_wfifo_we[1]~FF  (.D(\u_axi4_ctrl_0/n2656 ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), .Q(\u_axi4_ctrl_0/rc_wfifo_we[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/rc_wfifo_we[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_wfifo_we[2]~FF  (.D(\u_axi4_ctrl_0/n2661 ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), .Q(\u_axi4_ctrl_0/rc_wfifo_we[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/rc_wfifo_we[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_wfifo_we[3]~FF  (.D(\u_axi4_ctrl_0/n2666 ), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), .Q(\u_axi4_ctrl_0/rc_wfifo_we[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl_0/rc_wfifo_we[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_wfifo_we[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(515)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(515)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(508)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/w_wfifo_empty~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n71 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/w_wfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1106)
    defparam \u_axi4_ctrl_0/w_wfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_wfifo_empty~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_wfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_wfifo_empty~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_wfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/w_wfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/w_wfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n152 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n184 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n194 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n151 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n150 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n149 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n148 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n147 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n146 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n145 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n144 ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n183 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n182 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n181 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n180 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n179 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n178 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n177 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n176 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n193 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n192 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n191 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n190 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n189 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n188 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n187 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n186 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(n8651), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_axi4_ctrl_0/r_w_rst ), 
           .Q(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(508)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_cnt[2]~FF  (.D(\u_axi4_ctrl_0/n1073 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/n2551 ), .Q(\u_axi4_ctrl_0/rfifo_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(360)
    defparam \u_axi4_ctrl_0/rfifo_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[2]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_cnt[3]~FF  (.D(\u_axi4_ctrl_0/n1072 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/n2551 ), .Q(\u_axi4_ctrl_0/rfifo_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(360)
    defparam \u_axi4_ctrl_0/rfifo_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[3]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_cnt[4]~FF  (.D(\u_axi4_ctrl_0/n1071 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/n2551 ), .Q(\u_axi4_ctrl_0/rfifo_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(360)
    defparam \u_axi4_ctrl_0/rfifo_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[4]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/w_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(515)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/w_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(515)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/w_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(508)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/w_rfifo_empty~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n71 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/w_rfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1106)
    defparam \u_axi4_ctrl_0/w_rfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_rfifo_empty~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_rfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_rfifo_empty~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/w_rfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/w_rfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/w_rfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n152 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n184 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n194 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n151 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n150 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n149 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n148 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n147 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n146 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n145 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n144 ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1289)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n183 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n182 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n181 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n180 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n179 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n178 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n177 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n176 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n193 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n192 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n191 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n190 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n189 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n188 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n187 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n186 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1300)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1332)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1341)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1355)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1367)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[1][8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[1][8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(149)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/w_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(508)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF  (.D(\u_axi4_ctrl_0/n2677 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst_rclk ), 
           .Q(\u_axi4_ctrl_0/rc_rfifo_rd[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(427)
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF  (.D(\u_axi4_ctrl_0/n2682 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst_rclk ), 
           .Q(\u_axi4_ctrl_0/rc_rfifo_rd[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(427)
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rc_rfifo_rd[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[0]~FF  (.D(\u_axi4_ctrl_0/n1507 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[0]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[0]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[0]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[0]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[1]~FF  (.D(\u_axi4_ctrl_0/n1506 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[1]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[1]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[1]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[1]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[1]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[2]~FF  (.D(\u_axi4_ctrl_0/n1505 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[2]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[2]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[2]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[2]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[2]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[3]~FF  (.D(\u_axi4_ctrl_0/n1504 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[3]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[3]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[3]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[3]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[3]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[4]~FF  (.D(\u_axi4_ctrl_0/n1503 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[4]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[4]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[4]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[4]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[4]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[5]~FF  (.D(\u_axi4_ctrl_0/n1502 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[5]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[5]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[5]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[5]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[5]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[6]~FF  (.D(\u_axi4_ctrl_0/n1501 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[6]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[6]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[6]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[6]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[6]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[7]~FF  (.D(\u_axi4_ctrl_0/n1500 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[7]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[7]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[7]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[7]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[7]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[8]~FF  (.D(\u_axi4_ctrl_0/n1499 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[8]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[8]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[8]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[8]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[8]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[8]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[9]~FF  (.D(\u_axi4_ctrl_0/n1498 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[9]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[9]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[9]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[9]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[9]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[9]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[10]~FF  (.D(\u_axi4_ctrl_0/n1497 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[10]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[10]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[10]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[10]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[10]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[10]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[11]~FF  (.D(\u_axi4_ctrl_0/n1496 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[11]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[11]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[11]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[11]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[11]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[11]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[12]~FF  (.D(\u_axi4_ctrl_0/n1495 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[12]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[12]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[12]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[12]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[12]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[12]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[13]~FF  (.D(\u_axi4_ctrl_0/n1494 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[13]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[13]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[13]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[13]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[13]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[13]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[14]~FF  (.D(\u_axi4_ctrl_0/n1493 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[14]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[14]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[14]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[14]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[14]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[14]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_data[15]~FF  (.D(\u_axi4_ctrl_0/n1492 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_data[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \lcd_data[15]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_data[15]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_data[15]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_data[15]~FF .D_POLARITY = 1'b1;
    defparam \lcd_data[15]~FF .SR_SYNC = 1'b1;
    defparam \lcd_data[15]~FF .SR_VALUE = 1'b0;
    defparam \lcd_data[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF  (.D(\u_axi4_ctrl_0/n1491 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF  (.D(\u_axi4_ctrl_0/n1490 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF  (.D(\u_axi4_ctrl_0/n1489 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF  (.D(\u_axi4_ctrl_0/n1488 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF  (.D(\u_axi4_ctrl_0/n1487 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF  (.D(\u_axi4_ctrl_0/n1486 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF  (.D(\u_axi4_ctrl_0/n1485 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF  (.D(\u_axi4_ctrl_0/n1484 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF  (.D(\u_axi4_ctrl_0/n1483 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF  (.D(\u_axi4_ctrl_0/n1482 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF  (.D(\u_axi4_ctrl_0/n1481 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF  (.D(\u_axi4_ctrl_0/n1480 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF  (.D(\u_axi4_ctrl_0/n1479 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF  (.D(\u_axi4_ctrl_0/n1478 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF  (.D(\u_axi4_ctrl_0/n1477 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF  (.D(\u_axi4_ctrl_0/n1476 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF  (.D(\u_axi4_ctrl_0/n1475 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF  (.D(\u_axi4_ctrl_0/n1474 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF  (.D(\u_axi4_ctrl_0/n1473 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF  (.D(\u_axi4_ctrl_0/n1472 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF  (.D(\u_axi4_ctrl_0/n1471 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF  (.D(\u_axi4_ctrl_0/n1470 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF  (.D(\u_axi4_ctrl_0/n1469 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF  (.D(\u_axi4_ctrl_0/n1468 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF  (.D(\u_axi4_ctrl_0/n1467 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF  (.D(\u_axi4_ctrl_0/n1466 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF  (.D(\u_axi4_ctrl_0/n1465 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF  (.D(\u_axi4_ctrl_0/n1464 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF  (.D(\u_axi4_ctrl_0/n1463 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF  (.D(\u_axi4_ctrl_0/n1462 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF  (.D(\u_axi4_ctrl_0/n1461 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF  (.D(\u_axi4_ctrl_0/n1460 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF  (.D(\u_axi4_ctrl_0/n1459 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF  (.D(\u_axi4_ctrl_0/n1458 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF  (.D(\u_axi4_ctrl_0/n1457 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF  (.D(\u_axi4_ctrl_0/n1456 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF  (.D(\u_axi4_ctrl_0/n1455 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF  (.D(\u_axi4_ctrl_0/n1454 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF  (.D(\u_axi4_ctrl_0/n1453 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF  (.D(\u_axi4_ctrl_0/n1452 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF  (.D(\u_axi4_ctrl_0/n1451 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF  (.D(\u_axi4_ctrl_0/n1450 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF  (.D(\u_axi4_ctrl_0/n1449 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF  (.D(\u_axi4_ctrl_0/n1448 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF  (.D(\u_axi4_ctrl_0/n1447 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF  (.D(\u_axi4_ctrl_0/n1446 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF  (.D(\u_axi4_ctrl_0/n1445 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF  (.D(\u_axi4_ctrl_0/n1444 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF  (.D(\u_axi4_ctrl_0/n1443 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF  (.D(\u_axi4_ctrl_0/n1442 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF  (.D(\u_axi4_ctrl_0/n1441 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF  (.D(\u_axi4_ctrl_0/n1440 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF  (.D(\u_axi4_ctrl_0/n1439 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF  (.D(\u_axi4_ctrl_0/n1438 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF  (.D(\u_axi4_ctrl_0/n1437 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF  (.D(\u_axi4_ctrl_0/n1436 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF  (.D(\u_axi4_ctrl_0/n1435 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF  (.D(\u_axi4_ctrl_0/n1434 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF  (.D(\u_axi4_ctrl_0/n1433 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF  (.D(\u_axi4_ctrl_0/n1432 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF  (.D(\u_axi4_ctrl_0/n1431 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF  (.D(\u_axi4_ctrl_0/n1430 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF  (.D(\u_axi4_ctrl_0/n1429 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF  (.D(\u_axi4_ctrl_0/n1428 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF  (.D(\u_axi4_ctrl_0/n1427 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF  (.D(\u_axi4_ctrl_0/n1426 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF  (.D(\u_axi4_ctrl_0/n1425 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF  (.D(\u_axi4_ctrl_0/n1424 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF  (.D(\u_axi4_ctrl_0/n1423 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF  (.D(\u_axi4_ctrl_0/n1422 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF  (.D(\u_axi4_ctrl_0/n1421 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF  (.D(\u_axi4_ctrl_0/n1420 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF  (.D(\u_axi4_ctrl_0/n1419 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF  (.D(\u_axi4_ctrl_0/n1418 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF  (.D(\u_axi4_ctrl_0/n1417 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF  (.D(\u_axi4_ctrl_0/n1416 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF  (.D(\u_axi4_ctrl_0/n1415 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF  (.D(\u_axi4_ctrl_0/n1414 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF  (.D(\u_axi4_ctrl_0/n1413 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF  (.D(\u_axi4_ctrl_0/n1412 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF  (.D(\u_axi4_ctrl_0/n1411 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF  (.D(\u_axi4_ctrl_0/n1410 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF  (.D(\u_axi4_ctrl_0/n1409 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF  (.D(\u_axi4_ctrl_0/n1408 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF  (.D(\u_axi4_ctrl_0/n1407 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF  (.D(\u_axi4_ctrl_0/n1406 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF  (.D(\u_axi4_ctrl_0/n1405 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF  (.D(\u_axi4_ctrl_0/n1404 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF  (.D(\u_axi4_ctrl_0/n1403 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF  (.D(\u_axi4_ctrl_0/n1402 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF  (.D(\u_axi4_ctrl_0/n1401 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF  (.D(\u_axi4_ctrl_0/n1400 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF  (.D(\u_axi4_ctrl_0/n1399 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF  (.D(\u_axi4_ctrl_0/n1398 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF  (.D(\u_axi4_ctrl_0/n1397 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF  (.D(\u_axi4_ctrl_0/n1396 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF  (.D(\u_axi4_ctrl_0/n1395 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF  (.D(\u_axi4_ctrl_0/n1394 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF  (.D(\u_axi4_ctrl_0/n1393 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF  (.D(\u_axi4_ctrl_0/n1392 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF  (.D(\u_axi4_ctrl_0/n1391 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF  (.D(\u_axi4_ctrl_0/n1390 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF  (.D(\u_axi4_ctrl_0/n1389 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF  (.D(\u_axi4_ctrl_0/n1388 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF  (.D(\u_axi4_ctrl_0/n1387 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF  (.D(\u_axi4_ctrl_0/n1386 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF  (.D(\u_axi4_ctrl_0/n1385 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF  (.D(\u_axi4_ctrl_0/n1384 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF  (.D(\u_axi4_ctrl_0/n1383 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF  (.D(\u_axi4_ctrl_0/n1382 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF  (.D(\u_axi4_ctrl_0/n1381 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF  (.D(\u_axi4_ctrl_0/n1380 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/r_rframe_data_gen[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(440)
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/r_rframe_data_gen[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[2] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[3] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[4] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[5] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[6] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[7] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[8] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[9] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[10] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[11] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[12] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[13] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF  (.D(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[14] ), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), 
           .Q(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(453)
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[8]~FF  (.D(\u_axi4_ctrl_0/n1774 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[8]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[8]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[8]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[8]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[8]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[9]~FF  (.D(\u_axi4_ctrl_0/n1773 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[9]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[9]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[9]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[9]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[9]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[10]~FF  (.D(\u_axi4_ctrl_0/n1772 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[10]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[10]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[10]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[10]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[10]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[11]~FF  (.D(\u_axi4_ctrl_0/n1771 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[11]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[11]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[11]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[11]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[11]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[12]~FF  (.D(\u_axi4_ctrl_0/n1770 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[12]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[12]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[12]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[12]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[12]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[13]~FF  (.D(\u_axi4_ctrl_0/n1769 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[13]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[13]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[13]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[13]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[13]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[14]~FF  (.D(\u_axi4_ctrl_0/n1768 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[14]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[14]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[14]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[14]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[14]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[15]~FF  (.D(\u_axi4_ctrl_0/n1767 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[15]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[15]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[15]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[15]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[15]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[16]~FF  (.D(\u_axi4_ctrl_0/n1766 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[16]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[16]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[16]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[16]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[16]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[17]~FF  (.D(\u_axi4_ctrl_0/n1765 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[17]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[17]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[17]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[17]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[17]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[18]~FF  (.D(\u_axi4_ctrl_0/n1764 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[18]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[18]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[18]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[18]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[18]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[19]~FF  (.D(\u_axi4_ctrl_0/n1763 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[19]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[19]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[19]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[19]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[19]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[20]~FF  (.D(\u_axi4_ctrl_0/n1762 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[20]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[20]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[20]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[20]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[20]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ARADDR_0[21]~FF  (.D(\u_axi4_ctrl_0/n1761 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\u_axi4_ctrl_0/r_rfifo_rst ), .Q(\DdrCtrl_ARADDR_0[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(566)
    defparam \DdrCtrl_ARADDR_0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[21]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[21]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[21]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ARADDR_0[21]~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_ARADDR_0[21]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ARADDR_0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[4]~FF  (.D(DdrCtrl_RDATA_0[4]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[5]~FF  (.D(DdrCtrl_RDATA_0[5]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[6]~FF  (.D(DdrCtrl_RDATA_0[6]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[7]~FF  (.D(DdrCtrl_RDATA_0[7]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[8]~FF  (.D(DdrCtrl_RDATA_0[8]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[9]~FF  (.D(DdrCtrl_RDATA_0[9]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[10]~FF  (.D(DdrCtrl_RDATA_0[10]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[11]~FF  (.D(DdrCtrl_RDATA_0[11]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[12]~FF  (.D(DdrCtrl_RDATA_0[12]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[13]~FF  (.D(DdrCtrl_RDATA_0[13]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[14]~FF  (.D(DdrCtrl_RDATA_0[14]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[15]~FF  (.D(DdrCtrl_RDATA_0[15]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[16]~FF  (.D(DdrCtrl_RDATA_0[16]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[17]~FF  (.D(DdrCtrl_RDATA_0[17]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[18]~FF  (.D(DdrCtrl_RDATA_0[18]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[19]~FF  (.D(DdrCtrl_RDATA_0[19]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[20]~FF  (.D(DdrCtrl_RDATA_0[20]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[21]~FF  (.D(DdrCtrl_RDATA_0[21]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[22]~FF  (.D(DdrCtrl_RDATA_0[22]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[23]~FF  (.D(DdrCtrl_RDATA_0[23]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[24]~FF  (.D(DdrCtrl_RDATA_0[24]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[24]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[24]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[24]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[25]~FF  (.D(DdrCtrl_RDATA_0[25]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[25]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[25]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[25]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[26]~FF  (.D(DdrCtrl_RDATA_0[26]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[26]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[26]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[26]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[27]~FF  (.D(DdrCtrl_RDATA_0[27]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[27]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[27]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[27]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[28]~FF  (.D(DdrCtrl_RDATA_0[28]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[28]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[28]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[28]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[28]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[29]~FF  (.D(DdrCtrl_RDATA_0[29]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[29]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[29]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[29]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[29]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[30]~FF  (.D(DdrCtrl_RDATA_0[30]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[30]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[30]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[30]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[30]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[31]~FF  (.D(DdrCtrl_RDATA_0[31]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[31]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[31]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[31]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[31]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[32]~FF  (.D(DdrCtrl_RDATA_0[32]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[32]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[32]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[32]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[32]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[32]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[32]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[33]~FF  (.D(DdrCtrl_RDATA_0[33]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[33]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[33]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[33]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[33]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[33]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[33]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[34]~FF  (.D(DdrCtrl_RDATA_0[34]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[34]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[34]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[34]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[34]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[34]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[34]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[35]~FF  (.D(DdrCtrl_RDATA_0[35]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[35]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[35]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[35]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[35]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[35]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[35]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[36]~FF  (.D(DdrCtrl_RDATA_0[36]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[36]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[36]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[36]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[36]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[36]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[36]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[37]~FF  (.D(DdrCtrl_RDATA_0[37]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[37]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[37]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[37]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[37]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[37]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[37]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[38]~FF  (.D(DdrCtrl_RDATA_0[38]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[38]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[38]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[38]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[38]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[38]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[38]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[39]~FF  (.D(DdrCtrl_RDATA_0[39]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[39]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[39]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[39]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[39]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[39]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[39]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[40]~FF  (.D(DdrCtrl_RDATA_0[40]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[40]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[40]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[40]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[40]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[40]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[40]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[41]~FF  (.D(DdrCtrl_RDATA_0[41]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[41]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[41]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[41]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[41]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[41]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[41]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[42]~FF  (.D(DdrCtrl_RDATA_0[42]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[42]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[42]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[42]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[42]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[42]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[42]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[43]~FF  (.D(DdrCtrl_RDATA_0[43]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[43]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[43]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[43]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[43]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[43]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[43]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[44]~FF  (.D(DdrCtrl_RDATA_0[44]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[44]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[44]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[44]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[44]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[44]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[44]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[45]~FF  (.D(DdrCtrl_RDATA_0[45]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[45]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[45]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[45]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[45]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[45]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[45]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[46]~FF  (.D(DdrCtrl_RDATA_0[46]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[46]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[46]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[46]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[46]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[46]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[46]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[47]~FF  (.D(DdrCtrl_RDATA_0[47]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[47]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[47]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[47]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[47]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[47]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[47]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[48]~FF  (.D(DdrCtrl_RDATA_0[48]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[48]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[48]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[48]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[48]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[48]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[48]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[49]~FF  (.D(DdrCtrl_RDATA_0[49]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[49]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[49]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[49]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[49]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[49]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[49]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[50]~FF  (.D(DdrCtrl_RDATA_0[50]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[50]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[50]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[50]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[50]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[50]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[50]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[51]~FF  (.D(DdrCtrl_RDATA_0[51]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[51]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[51]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[51]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[51]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[51]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[51]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[52]~FF  (.D(DdrCtrl_RDATA_0[52]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[52]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[52]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[52]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[52]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[52]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[52]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[53]~FF  (.D(DdrCtrl_RDATA_0[53]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[53]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[53]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[53]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[53]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[53]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[53]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[54]~FF  (.D(DdrCtrl_RDATA_0[54]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[54]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[54]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[54]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[54]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[54]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[54]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[55]~FF  (.D(DdrCtrl_RDATA_0[55]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[55]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[55]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[55]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[55]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[55]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[55]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[56]~FF  (.D(DdrCtrl_RDATA_0[56]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[56]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[56]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[56]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[56]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[56]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[56]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[57]~FF  (.D(DdrCtrl_RDATA_0[57]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[57]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[57]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[57]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[57]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[57]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[57]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[58]~FF  (.D(DdrCtrl_RDATA_0[58]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[58]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[58]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[58]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[58]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[58]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[58]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[59]~FF  (.D(DdrCtrl_RDATA_0[59]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[59]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[59]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[59]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[59]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[59]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[59]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[60]~FF  (.D(DdrCtrl_RDATA_0[60]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[60]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[60]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[60]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[60]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[60]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[60]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[61]~FF  (.D(DdrCtrl_RDATA_0[61]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[61]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[61]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[61]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[61]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[61]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[61]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[62]~FF  (.D(DdrCtrl_RDATA_0[62]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[62]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[62]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[62]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[62]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[62]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[62]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[63]~FF  (.D(DdrCtrl_RDATA_0[63]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[63]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[63]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[63]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[63]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[63]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[63]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[64]~FF  (.D(DdrCtrl_RDATA_0[64]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[64]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[64]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[64]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[64]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[64]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[64]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[65]~FF  (.D(DdrCtrl_RDATA_0[65]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[65]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[65]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[65]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[65]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[65]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[65]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[66]~FF  (.D(DdrCtrl_RDATA_0[66]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[66]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[66]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[66]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[66]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[66]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[66]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[67]~FF  (.D(DdrCtrl_RDATA_0[67]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[67]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[67]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[67]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[67]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[67]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[67]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[68]~FF  (.D(DdrCtrl_RDATA_0[68]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[68]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[68]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[68]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[68]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[68]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[68]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[69]~FF  (.D(DdrCtrl_RDATA_0[69]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[69]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[69]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[69]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[69]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[69]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[69]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[70]~FF  (.D(DdrCtrl_RDATA_0[70]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[70]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[70]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[70]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[70]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[70]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[70]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[71]~FF  (.D(DdrCtrl_RDATA_0[71]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[71]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[71]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[71]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[71]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[71]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[71]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[72]~FF  (.D(DdrCtrl_RDATA_0[72]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[72]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[72]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[72]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[72]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[72]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[72]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[73]~FF  (.D(DdrCtrl_RDATA_0[73]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[73]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[73]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[73]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[73]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[73]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[73]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[74]~FF  (.D(DdrCtrl_RDATA_0[74]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[74]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[74]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[74]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[74]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[74]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[74]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[75]~FF  (.D(DdrCtrl_RDATA_0[75]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[75]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[75]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[75]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[75]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[75]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[75]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[76]~FF  (.D(DdrCtrl_RDATA_0[76]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[76]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[76]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[76]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[76]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[76]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[76]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[77]~FF  (.D(DdrCtrl_RDATA_0[77]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[77]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[77]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[77]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[77]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[77]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[77]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[78]~FF  (.D(DdrCtrl_RDATA_0[78]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[78]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[78]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[78]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[78]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[78]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[78]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[79]~FF  (.D(DdrCtrl_RDATA_0[79]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[79]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[79]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[79]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[79]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[79]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[79]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[80]~FF  (.D(DdrCtrl_RDATA_0[80]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[80]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[80]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[80]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[80]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[80]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[80]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[81]~FF  (.D(DdrCtrl_RDATA_0[81]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[81]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[81]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[81]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[81]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[81]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[81]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[82]~FF  (.D(DdrCtrl_RDATA_0[82]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[82]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[82]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[82]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[82]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[82]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[82]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[83]~FF  (.D(DdrCtrl_RDATA_0[83]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[83]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[83]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[83]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[83]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[83]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[83]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[84]~FF  (.D(DdrCtrl_RDATA_0[84]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[84]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[84]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[84]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[84]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[84]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[84]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[85]~FF  (.D(DdrCtrl_RDATA_0[85]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[85]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[85]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[85]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[85]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[85]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[85]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[86]~FF  (.D(DdrCtrl_RDATA_0[86]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[86]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[86]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[86]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[86]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[86]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[86]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[87]~FF  (.D(DdrCtrl_RDATA_0[87]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[87]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[87]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[87]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[87]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[87]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[87]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[88]~FF  (.D(DdrCtrl_RDATA_0[88]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[88]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[88]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[88]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[88]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[88]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[88]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[89]~FF  (.D(DdrCtrl_RDATA_0[89]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[89]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[89]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[89]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[89]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[89]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[89]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[90]~FF  (.D(DdrCtrl_RDATA_0[90]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[90]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[90]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[90]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[90]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[90]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[90]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[91]~FF  (.D(DdrCtrl_RDATA_0[91]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[91]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[91]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[91]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[91]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[91]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[91]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[92]~FF  (.D(DdrCtrl_RDATA_0[92]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[92]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[92]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[92]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[92]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[92]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[92]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[93]~FF  (.D(DdrCtrl_RDATA_0[93]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[93]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[93]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[93]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[93]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[93]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[93]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[94]~FF  (.D(DdrCtrl_RDATA_0[94]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[94]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[94]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[94]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[94]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[94]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[94]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[95]~FF  (.D(DdrCtrl_RDATA_0[95]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[95]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[95]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[95]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[95]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[95]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[95]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[96]~FF  (.D(DdrCtrl_RDATA_0[96]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[96]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[96]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[96]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[96]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[96]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[96]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[97]~FF  (.D(DdrCtrl_RDATA_0[97]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[97]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[97]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[97]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[97]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[97]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[97]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[98]~FF  (.D(DdrCtrl_RDATA_0[98]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[98]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[98]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[98]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[98]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[98]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[98]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[99]~FF  (.D(DdrCtrl_RDATA_0[99]), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[99]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[99]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[99]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[99]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[99]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[99]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[100]~FF  (.D(DdrCtrl_RDATA_0[100]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[100]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[100]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[100]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[100]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[100]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[100]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[101]~FF  (.D(DdrCtrl_RDATA_0[101]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[101]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[101]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[101]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[101]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[101]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[101]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[102]~FF  (.D(DdrCtrl_RDATA_0[102]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[102]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[102]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[102]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[102]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[102]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[102]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[103]~FF  (.D(DdrCtrl_RDATA_0[103]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[103]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[103]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[103]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[103]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[103]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[103]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[104]~FF  (.D(DdrCtrl_RDATA_0[104]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[104]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[104]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[104]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[104]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[104]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[104]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[105]~FF  (.D(DdrCtrl_RDATA_0[105]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[105]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[105]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[105]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[105]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[105]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[105]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[106]~FF  (.D(DdrCtrl_RDATA_0[106]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[106]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[106]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[106]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[106]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[106]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[106]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[107]~FF  (.D(DdrCtrl_RDATA_0[107]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[107]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[107]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[107]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[107]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[107]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[107]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[108]~FF  (.D(DdrCtrl_RDATA_0[108]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[108]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[108]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[108]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[108]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[108]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[108]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[109]~FF  (.D(DdrCtrl_RDATA_0[109]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[109]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[109]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[109]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[109]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[109]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[109]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[110]~FF  (.D(DdrCtrl_RDATA_0[110]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[110]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[110]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[110]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[110]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[110]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[110]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[111]~FF  (.D(DdrCtrl_RDATA_0[111]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[111]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[111]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[111]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[111]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[111]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[111]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[112]~FF  (.D(DdrCtrl_RDATA_0[112]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[112]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[112]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[112]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[112]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[112]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[112]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[113]~FF  (.D(DdrCtrl_RDATA_0[113]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[113]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[113]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[113]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[113]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[113]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[113]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[114]~FF  (.D(DdrCtrl_RDATA_0[114]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[114]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[114]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[114]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[114]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[114]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[114]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[115]~FF  (.D(DdrCtrl_RDATA_0[115]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[115]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[115]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[115]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[115]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[115]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[115]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[116]~FF  (.D(DdrCtrl_RDATA_0[116]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[116]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[116]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[116]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[116]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[116]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[116]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[117]~FF  (.D(DdrCtrl_RDATA_0[117]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[117]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[117]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[117]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[117]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[117]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[117]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[118]~FF  (.D(DdrCtrl_RDATA_0[118]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[118]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[118]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[118]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[118]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[118]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[118]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[119]~FF  (.D(DdrCtrl_RDATA_0[119]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[119]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[119]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[119]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[119]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[119]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[119]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[120]~FF  (.D(DdrCtrl_RDATA_0[120]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[120]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[120]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[120]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[120]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[120]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[120]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[121]~FF  (.D(DdrCtrl_RDATA_0[121]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[121]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[121]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[121]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[121]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[121]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[121]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[122]~FF  (.D(DdrCtrl_RDATA_0[122]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[122]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[122]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[122]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[122]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[122]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[122]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[123]~FF  (.D(DdrCtrl_RDATA_0[123]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[123]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[123]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[123]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[123]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[123]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[123]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[124]~FF  (.D(DdrCtrl_RDATA_0[124]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[124]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[124]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[124]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[124]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[124]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[124]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[125]~FF  (.D(DdrCtrl_RDATA_0[125]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[125]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[125]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[125]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[125]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[125]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[125]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[126]~FF  (.D(DdrCtrl_RDATA_0[126]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[126]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[126]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[126]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[126]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[126]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[126]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl_0/rfifo_wdata[127]~FF  (.D(DdrCtrl_RDATA_0[127]), 
           .CE(1'b1), .CLK(\Axi0Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl_0/rfifo_wdata[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(610)
    defparam \u_axi4_ctrl_0/rfifo_wdata[127]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[127]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[127]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[127]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[127]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl_0/rfifo_wdata[127]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl_0/rfifo_wdata[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AWADDR_0[23]~FF  (.D(\u_axi4_ctrl_0/n2772 ), .CE(1'b1), 
           .CLK(\Axi0Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\DdrCtrl_AWADDR_0[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(154)
    defparam \DdrCtrl_AWADDR_0[23]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[23]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[23]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AWADDR_0[23]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AWADDR_0[23]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AWADDR_0[23]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AWADDR_0[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[0]~FF  (.D(\u_lcd_driver/n96 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_hs~FF  (.D(\u_lcd_driver/n51 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_hs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \lcd_hs~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_hs~FF .CE_POLARITY = 1'b1;
    defparam \lcd_hs~FF .SR_POLARITY = 1'b1;
    defparam \lcd_hs~FF .D_POLARITY = 1'b1;
    defparam \lcd_hs~FF .SR_SYNC = 1'b1;
    defparam \lcd_hs~FF .SR_VALUE = 1'b0;
    defparam \lcd_hs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_vs~FF  (.D(\u_lcd_driver/n113 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_vs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \lcd_vs~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_vs~FF .CE_POLARITY = 1'b1;
    defparam \lcd_vs~FF .SR_POLARITY = 1'b1;
    defparam \lcd_vs~FF .D_POLARITY = 1'b1;
    defparam \lcd_vs~FF .SR_SYNC = 1'b1;
    defparam \lcd_vs~FF .SR_VALUE = 1'b0;
    defparam \lcd_vs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_dv~FF  (.D(\u_lcd_driver/n125 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_dv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_dv~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_request~FF  (.D(\u_lcd_driver/n194 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_request)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_request~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_request~FF .CE_POLARITY = 1'b1;
    defparam \lcd_request~FF .SR_POLARITY = 1'b1;
    defparam \lcd_request~FF .D_POLARITY = 1'b1;
    defparam \lcd_request~FF .SR_SYNC = 1'b1;
    defparam \lcd_request~FF .SR_VALUE = 1'b0;
    defparam \lcd_request~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[0]~FF  (.D(\u_lcd_driver/hcnt[0] ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[0]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[0]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[0]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[0]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[0]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[0]~FF  (.D(n1662), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[0]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[0]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[0]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[0]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[0]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[0]~FF  (.D(\u_lcd_driver/n34 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[1]~FF  (.D(\u_lcd_driver/n95 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[2]~FF  (.D(\u_lcd_driver/n94 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[3]~FF  (.D(\u_lcd_driver/n93 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[4]~FF  (.D(\u_lcd_driver/n92 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[5]~FF  (.D(\u_lcd_driver/n91 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[6]~FF  (.D(\u_lcd_driver/n90 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[7]~FF  (.D(\u_lcd_driver/n89 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[8]~FF  (.D(\u_lcd_driver/n88 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[9]~FF  (.D(\u_lcd_driver/n87 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[10]~FF  (.D(\u_lcd_driver/n86 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[11]~FF  (.D(\u_lcd_driver/n85 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[23]~FF  (.D(n733), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[23]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[23]~FF .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[23]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[1]~FF  (.D(n1657), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[1]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[1]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[1]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[1]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[1]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[2]~FF  (.D(n4173), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[2]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[2]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[2]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[2]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[2]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[3]~FF  (.D(n4171), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[3]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[3]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[3]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[3]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[3]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[4]~FF  (.D(n4169), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[4]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[4]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[4]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[4]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[4]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[5]~FF  (.D(n4167), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[5]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[5]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[5]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[5]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[5]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[6]~FF  (.D(n4165), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[6]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[6]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[6]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[6]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[6]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[7]~FF  (.D(n4163), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[7]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[7]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[7]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[7]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[7]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[8]~FF  (.D(n4161), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[8]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[8]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[8]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[8]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[8]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[9]~FF  (.D(n4159), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[9]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[9]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[9]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[9]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[9]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[10]~FF  (.D(n4157), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[10]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[10]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[10]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[10]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[10]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_xpos[11]~FF  (.D(n4156), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_xpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_xpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_xpos[11]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_xpos[11]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_xpos[11]~FF .D_POLARITY = 1'b1;
    defparam \lcd_xpos[11]~FF .SR_SYNC = 1'b1;
    defparam \lcd_xpos[11]~FF .SR_VALUE = 1'b0;
    defparam \lcd_xpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[1]~FF  (.D(n4154), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[1]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[1]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[1]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[1]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[1]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[2]~FF  (.D(n4152), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[2]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[2]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[2]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[2]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[2]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[3]~FF  (.D(n4150), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[3]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[3]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[3]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[3]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[3]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[4]~FF  (.D(n4148), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[4]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[4]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[4]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[4]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[4]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[5]~FF  (.D(n4146), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[5]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[5]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[5]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[5]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[5]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[6]~FF  (.D(n4144), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[6]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[6]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[6]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[6]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[6]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[7]~FF  (.D(n4142), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[7]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[7]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[7]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[7]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[7]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[8]~FF  (.D(n4140), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[8]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[8]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[8]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[8]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[8]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[9]~FF  (.D(n4138), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[9]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[9]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[9]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[9]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[9]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[10]~FF  (.D(n4136), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[10]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[10]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[10]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[10]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[10]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_ypos[11]~FF  (.D(n4135), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\lcd_ypos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(149)
    defparam \lcd_ypos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_ypos[11]~FF .CE_POLARITY = 1'b1;
    defparam \lcd_ypos[11]~FF .SR_POLARITY = 1'b1;
    defparam \lcd_ypos[11]~FF .D_POLARITY = 1'b1;
    defparam \lcd_ypos[11]~FF .SR_SYNC = 1'b1;
    defparam \lcd_ypos[11]~FF .SR_VALUE = 1'b0;
    defparam \lcd_ypos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[1]~FF  (.D(\u_lcd_driver/n33 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[2]~FF  (.D(\u_lcd_driver/n32 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[3]~FF  (.D(\u_lcd_driver/n31 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[4]~FF  (.D(\u_lcd_driver/n30 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[5]~FF  (.D(\u_lcd_driver/n29 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[6]~FF  (.D(\u_lcd_driver/n28 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[7]~FF  (.D(\u_lcd_driver/n27 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[8]~FF  (.D(\u_lcd_driver/n26 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[9]~FF  (.D(\u_lcd_driver/n25 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[10]~FF  (.D(\u_lcd_driver/n24 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[11]~FF  (.D(\u_lcd_driver/n23 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[0]~FF  (.D(\u_black_pixel_avg/n175 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[0]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[0]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[0]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[0]~FF  (.D(\u_black_pixel_avg/n208 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[0]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[0]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[0]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[1]~FF  (.D(\u_black_pixel_avg/n141 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[1]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[1]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[1]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[0]~FF  (.D(\u_black_pixel_avg/n142 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[0]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[0]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[0]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[1]~FF  (.D(\u_black_pixel_avg/n174 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[1]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[1]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[1]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[2]~FF  (.D(\u_black_pixel_avg/n173 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[2]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[2]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[2]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[3]~FF  (.D(\u_black_pixel_avg/n172 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[3]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[3]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[3]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[4]~FF  (.D(\u_black_pixel_avg/n171 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[4]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[4]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[4]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[5]~FF  (.D(\u_black_pixel_avg/n170 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[5]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[5]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[5]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[6]~FF  (.D(\u_black_pixel_avg/n169 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[6]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[6]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[6]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[7]~FF  (.D(\u_black_pixel_avg/n168 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[7]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[7]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[7]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[8]~FF  (.D(\u_black_pixel_avg/n167 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[8]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[8]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[8]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[9]~FF  (.D(\u_black_pixel_avg/n166 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[9]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[9]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[9]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[10]~FF  (.D(\u_black_pixel_avg/n165 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[10]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[10]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[10]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[11]~FF  (.D(\u_black_pixel_avg/n164 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[11]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[11]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[11]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[12]~FF  (.D(\u_black_pixel_avg/n163 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[12]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[12]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[12]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[13]~FF  (.D(\u_black_pixel_avg/n162 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[13]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[13]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[13]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[14]~FF  (.D(\u_black_pixel_avg/n161 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[14]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[14]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[14]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[15]~FF  (.D(\u_black_pixel_avg/n160 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[15]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[15]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[15]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[16]~FF  (.D(\u_black_pixel_avg/n159 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[16]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[16]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[16]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[17]~FF  (.D(\u_black_pixel_avg/n158 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[17]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[17]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[17]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[18]~FF  (.D(\u_black_pixel_avg/n157 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[18]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[18]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[18]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[19]~FF  (.D(\u_black_pixel_avg/n156 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[19]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[19]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[19]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[20]~FF  (.D(\u_black_pixel_avg/n155 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[20]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[20]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[20]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[20]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[21]~FF  (.D(\u_black_pixel_avg/n154 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[21]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[21]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[21]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[21]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[22]~FF  (.D(\u_black_pixel_avg/n153 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[22]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[22]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[22]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[22]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[23]~FF  (.D(\u_black_pixel_avg/n152 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[23]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[23]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[23]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[23]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[24]~FF  (.D(\u_black_pixel_avg/n151 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[24]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[24]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[24]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[24]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[25]~FF  (.D(\u_black_pixel_avg/n150 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[25]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[25]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[25]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[25]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[26]~FF  (.D(\u_black_pixel_avg/n149 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[26]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[26]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[26]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[26]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[27]~FF  (.D(\u_black_pixel_avg/n148 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[27]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[27]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[27]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[27]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[28]~FF  (.D(\u_black_pixel_avg/n147 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[28]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[28]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[28]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[28]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[29]~FF  (.D(\u_black_pixel_avg/n146 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[29]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[29]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[29]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[29]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[30]~FF  (.D(\u_black_pixel_avg/n145 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[30]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[30]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[30]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[30]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/y_sum[31]~FF  (.D(\u_black_pixel_avg/n144 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/y_sum[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/y_sum[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[31]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/y_sum[31]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/y_sum[31]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/y_sum[31]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/y_sum[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[1]~FF  (.D(\u_black_pixel_avg/n207 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[1]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[1]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[1]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[2]~FF  (.D(\u_black_pixel_avg/n206 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[2]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[2]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[2]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[3]~FF  (.D(\u_black_pixel_avg/n205 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[3]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[3]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[3]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[4]~FF  (.D(\u_black_pixel_avg/n204 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[4]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[4]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[4]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[5]~FF  (.D(\u_black_pixel_avg/n203 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[5]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[5]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[5]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[6]~FF  (.D(\u_black_pixel_avg/n202 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[6]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[6]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[6]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[7]~FF  (.D(\u_black_pixel_avg/n201 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[7]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[7]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[7]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[8]~FF  (.D(\u_black_pixel_avg/n200 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[8]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[8]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[8]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[9]~FF  (.D(\u_black_pixel_avg/n199 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[9]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[9]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[9]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[10]~FF  (.D(\u_black_pixel_avg/n198 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[10]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[10]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[10]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[11]~FF  (.D(\u_black_pixel_avg/n197 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[11]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[11]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[11]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[12]~FF  (.D(\u_black_pixel_avg/n196 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[12]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[12]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[12]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[13]~FF  (.D(\u_black_pixel_avg/n195 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[13]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[13]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[13]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[14]~FF  (.D(\u_black_pixel_avg/n194 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[14]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[14]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[14]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[15]~FF  (.D(\u_black_pixel_avg/n193 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[15]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[15]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[15]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[16]~FF  (.D(\u_black_pixel_avg/n192 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[16]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[16]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[16]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[17]~FF  (.D(\u_black_pixel_avg/n191 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[17]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[17]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[17]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[18]~FF  (.D(\u_black_pixel_avg/n190 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[18]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[18]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[18]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[19]~FF  (.D(\u_black_pixel_avg/n189 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[19]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[19]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[19]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[20]~FF  (.D(\u_black_pixel_avg/n188 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[20]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[20]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[20]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[20]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[21]~FF  (.D(\u_black_pixel_avg/n187 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[21]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[21]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[21]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[21]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[22]~FF  (.D(\u_black_pixel_avg/n186 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[22]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[22]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[22]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[22]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[23]~FF  (.D(\u_black_pixel_avg/n185 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[23]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[23]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[23]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[23]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[24]~FF  (.D(\u_black_pixel_avg/n184 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[24]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[24]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[24]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[24]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[25]~FF  (.D(\u_black_pixel_avg/n183 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[25]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[25]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[25]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[25]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[26]~FF  (.D(\u_black_pixel_avg/n182 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[26]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[26]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[26]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[26]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[27]~FF  (.D(\u_black_pixel_avg/n181 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[27]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[27]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[27]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[27]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[28]~FF  (.D(\u_black_pixel_avg/n180 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[28]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[28]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[28]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[28]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[29]~FF  (.D(\u_black_pixel_avg/n179 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[29]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[29]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[29]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[29]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[30]~FF  (.D(\u_black_pixel_avg/n178 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[30]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[30]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[30]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[30]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/black_pixel_count[31]~FF  (.D(\u_black_pixel_avg/n177 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/black_pixel_count[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/black_pixel_count[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[31]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[31]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[31]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/black_pixel_count[31]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/black_pixel_count[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \x_avg_black[6]~FF  (.D(\u_black_pixel_avg/n483 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\x_avg_black[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \x_avg_black[6]~FF .CLK_POLARITY = 1'b1;
    defparam \x_avg_black[6]~FF .CE_POLARITY = 1'b1;
    defparam \x_avg_black[6]~FF .SR_POLARITY = 1'b1;
    defparam \x_avg_black[6]~FF .D_POLARITY = 1'b1;
    defparam \x_avg_black[6]~FF .SR_SYNC = 1'b1;
    defparam \x_avg_black[6]~FF .SR_VALUE = 1'b0;
    defparam \x_avg_black[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \x_avg_black[7]~FF  (.D(\u_black_pixel_avg/n482 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\x_avg_black[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \x_avg_black[7]~FF .CLK_POLARITY = 1'b1;
    defparam \x_avg_black[7]~FF .CE_POLARITY = 1'b1;
    defparam \x_avg_black[7]~FF .SR_POLARITY = 1'b1;
    defparam \x_avg_black[7]~FF .D_POLARITY = 1'b1;
    defparam \x_avg_black[7]~FF .SR_SYNC = 1'b1;
    defparam \x_avg_black[7]~FF .SR_VALUE = 1'b0;
    defparam \x_avg_black[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \x_avg_black[8]~FF  (.D(\u_black_pixel_avg/n481 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\x_avg_black[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \x_avg_black[8]~FF .CLK_POLARITY = 1'b1;
    defparam \x_avg_black[8]~FF .CE_POLARITY = 1'b1;
    defparam \x_avg_black[8]~FF .SR_POLARITY = 1'b1;
    defparam \x_avg_black[8]~FF .D_POLARITY = 1'b1;
    defparam \x_avg_black[8]~FF .SR_SYNC = 1'b1;
    defparam \x_avg_black[8]~FF .SR_VALUE = 1'b0;
    defparam \x_avg_black[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \x_avg_black[9]~FF  (.D(\u_black_pixel_avg/n480 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\x_avg_black[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \x_avg_black[9]~FF .CLK_POLARITY = 1'b1;
    defparam \x_avg_black[9]~FF .CE_POLARITY = 1'b1;
    defparam \x_avg_black[9]~FF .SR_POLARITY = 1'b1;
    defparam \x_avg_black[9]~FF .D_POLARITY = 1'b1;
    defparam \x_avg_black[9]~FF .SR_SYNC = 1'b1;
    defparam \x_avg_black[9]~FF .SR_VALUE = 1'b0;
    defparam \x_avg_black[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \x_avg_black[10]~FF  (.D(\u_black_pixel_avg/n479 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\x_avg_black[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \x_avg_black[10]~FF .CLK_POLARITY = 1'b1;
    defparam \x_avg_black[10]~FF .CE_POLARITY = 1'b1;
    defparam \x_avg_black[10]~FF .SR_POLARITY = 1'b1;
    defparam \x_avg_black[10]~FF .D_POLARITY = 1'b1;
    defparam \x_avg_black[10]~FF .SR_SYNC = 1'b1;
    defparam \x_avg_black[10]~FF .SR_VALUE = 1'b0;
    defparam \x_avg_black[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \x_avg_black[11]~FF  (.D(\u_black_pixel_avg/n478 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\x_avg_black[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \x_avg_black[11]~FF .CLK_POLARITY = 1'b1;
    defparam \x_avg_black[11]~FF .CE_POLARITY = 1'b1;
    defparam \x_avg_black[11]~FF .SR_POLARITY = 1'b1;
    defparam \x_avg_black[11]~FF .D_POLARITY = 1'b1;
    defparam \x_avg_black[11]~FF .SR_SYNC = 1'b1;
    defparam \x_avg_black[11]~FF .SR_VALUE = 1'b0;
    defparam \x_avg_black[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[3]~FF  (.D(\u_black_pixel_avg/n499 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[3]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[3]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[3]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[3]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[3]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[3]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[4]~FF  (.D(\u_black_pixel_avg/n498 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[4]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[4]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[4]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[4]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[4]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[4]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[5]~FF  (.D(\u_black_pixel_avg/n497 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[5]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[5]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[5]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[5]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[5]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[5]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[6]~FF  (.D(\u_black_pixel_avg/n496 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[6]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[6]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[6]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[6]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[6]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[6]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[7]~FF  (.D(\u_black_pixel_avg/n495 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[7]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[7]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[7]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[7]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[7]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[7]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[8]~FF  (.D(\u_black_pixel_avg/n494 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[8]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[8]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[8]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[8]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[8]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[8]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[9]~FF  (.D(\u_black_pixel_avg/n493 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[9]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[9]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[9]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[9]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[9]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[9]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[10]~FF  (.D(\u_black_pixel_avg/n492 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[10]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[10]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[10]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[10]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[10]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[10]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \y_avg_black[11]~FF  (.D(\u_black_pixel_avg/n491 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\y_avg_black[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(50)
    defparam \y_avg_black[11]~FF .CLK_POLARITY = 1'b1;
    defparam \y_avg_black[11]~FF .CE_POLARITY = 1'b1;
    defparam \y_avg_black[11]~FF .SR_POLARITY = 1'b1;
    defparam \y_avg_black[11]~FF .D_POLARITY = 1'b1;
    defparam \y_avg_black[11]~FF .SR_SYNC = 1'b1;
    defparam \y_avg_black[11]~FF .SR_VALUE = 1'b0;
    defparam \y_avg_black[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[2]~FF  (.D(\u_black_pixel_avg/n140 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[2]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[2]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[2]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[3]~FF  (.D(\u_black_pixel_avg/n139 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[3]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[3]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[3]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[4]~FF  (.D(\u_black_pixel_avg/n138 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[4]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[4]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[4]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[5]~FF  (.D(\u_black_pixel_avg/n137 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[5]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[5]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[5]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[6]~FF  (.D(\u_black_pixel_avg/n136 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[6]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[6]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[6]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[7]~FF  (.D(\u_black_pixel_avg/n135 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[7]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[7]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[7]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[8]~FF  (.D(\u_black_pixel_avg/n134 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[8]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[8]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[8]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[9]~FF  (.D(\u_black_pixel_avg/n133 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[9]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[9]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[9]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[10]~FF  (.D(\u_black_pixel_avg/n132 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[10]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[10]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[10]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[11]~FF  (.D(\u_black_pixel_avg/n131 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[11]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[11]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[11]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[12]~FF  (.D(\u_black_pixel_avg/n130 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[12]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[12]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[12]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[13]~FF  (.D(\u_black_pixel_avg/n129 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[13]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[13]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[13]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[14]~FF  (.D(\u_black_pixel_avg/n128 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[14]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[14]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[14]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[15]~FF  (.D(\u_black_pixel_avg/n127 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[15]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[15]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[15]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[16]~FF  (.D(\u_black_pixel_avg/n126 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[16]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[16]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[16]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[17]~FF  (.D(\u_black_pixel_avg/n125 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[17]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[17]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[17]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[18]~FF  (.D(\u_black_pixel_avg/n124 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[18]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[18]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[18]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[19]~FF  (.D(\u_black_pixel_avg/n123 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[19]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[19]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[19]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[20]~FF  (.D(\u_black_pixel_avg/n122 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[20]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[20]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[20]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[20]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[21]~FF  (.D(\u_black_pixel_avg/n121 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[21]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[21]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[21]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[21]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[22]~FF  (.D(\u_black_pixel_avg/n120 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[22]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[22]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[22]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[22]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[23]~FF  (.D(\u_black_pixel_avg/n119 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[23]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[23]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[23]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[23]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[24]~FF  (.D(\u_black_pixel_avg/n118 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[24]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[24]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[24]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[24]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[25]~FF  (.D(\u_black_pixel_avg/n117 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[25]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[25]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[25]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[25]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[26]~FF  (.D(\u_black_pixel_avg/n116 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[26]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[26]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[26]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[26]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[27]~FF  (.D(\u_black_pixel_avg/n115 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[27]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[27]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[27]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[27]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[28]~FF  (.D(\u_black_pixel_avg/n114 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[28]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[28]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[28]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[28]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[29]~FF  (.D(\u_black_pixel_avg/n113 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[29]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[29]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[29]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[29]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[30]~FF  (.D(\u_black_pixel_avg/n112 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[30]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[30]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[30]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[30]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_black_pixel_avg/x_sum[31]~FF  (.D(\u_black_pixel_avg/n111 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_vs), .Q(\u_black_pixel_avg/x_sum[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(41)
    defparam \u_black_pixel_avg/x_sum[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[31]~FF .SR_POLARITY = 1'b0;
    defparam \u_black_pixel_avg/x_sum[31]~FF .D_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/x_sum[31]~FF .SR_SYNC = 1'b1;
    defparam \u_black_pixel_avg/x_sum[31]~FF .SR_VALUE = 1'b0;
    defparam \u_black_pixel_avg/x_sum[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/key0_last~FF  (.D(key0), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\u_state_machine/key0_last )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(28)
    defparam \u_state_machine/key0_last~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/key0_last~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/key0_last~FF .SR_POLARITY = 1'b1;
    defparam \u_state_machine/key0_last~FF .D_POLARITY = 1'b0;
    defparam \u_state_machine/key0_last~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/key0_last~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/key0_last~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/current_state.WAITING~FF  (.D(\u_state_machine/next_state.WAITING ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_state_machine/current_state.WAITING )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/current_state.WAITING~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/current_state.WAITING~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/current_state.WAITING~FF .SR_POLARITY = 1'b1;
    defparam \u_state_machine/current_state.WAITING~FF .D_POLARITY = 1'b0;
    defparam \u_state_machine/current_state.WAITING~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/current_state.WAITING~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/current_state.WAITING~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[0]~FF  (.D(\u_state_machine/n113 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[0]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[0]~FF .D_POLARITY = 1'b1;
    defparam \led_data[0]~FF .SR_SYNC = 1'b1;
    defparam \led_data[0]~FF .SR_VALUE = 1'b0;
    defparam \led_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/current_state.WORKING~FF  (.D(\u_state_machine/next_state.WORKING ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_state_machine/current_state.WORKING )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/current_state.WORKING~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/current_state.WORKING~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/current_state.WORKING~FF .SR_POLARITY = 1'b1;
    defparam \u_state_machine/current_state.WORKING~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/current_state.WORKING~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/current_state.WORKING~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/current_state.WORKING~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[0]~FF  (.D(\u_state_machine/n99 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[0]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[0]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[0]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \zone_bit0~FF  (.D(\u_state_machine/n114 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(zone_bit0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \zone_bit0~FF .CLK_POLARITY = 1'b1;
    defparam \zone_bit0~FF .CE_POLARITY = 1'b1;
    defparam \zone_bit0~FF .SR_POLARITY = 1'b1;
    defparam \zone_bit0~FF .D_POLARITY = 1'b1;
    defparam \zone_bit0~FF .SR_SYNC = 1'b1;
    defparam \zone_bit0~FF .SR_VALUE = 1'b0;
    defparam \zone_bit0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \zone_bit1~FF  (.D(\u_state_machine/n115 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(zone_bit1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \zone_bit1~FF .CLK_POLARITY = 1'b1;
    defparam \zone_bit1~FF .CE_POLARITY = 1'b1;
    defparam \zone_bit1~FF .SR_POLARITY = 1'b1;
    defparam \zone_bit1~FF .D_POLARITY = 1'b1;
    defparam \zone_bit1~FF .SR_SYNC = 1'b1;
    defparam \zone_bit1~FF .SR_VALUE = 1'b0;
    defparam \zone_bit1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \zone_bit2~FF  (.D(\u_state_machine/n116 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(zone_bit2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \zone_bit2~FF .CLK_POLARITY = 1'b1;
    defparam \zone_bit2~FF .CE_POLARITY = 1'b1;
    defparam \zone_bit2~FF .SR_POLARITY = 1'b1;
    defparam \zone_bit2~FF .D_POLARITY = 1'b1;
    defparam \zone_bit2~FF .SR_SYNC = 1'b1;
    defparam \zone_bit2~FF .SR_VALUE = 1'b0;
    defparam \zone_bit2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/next_state.WAITING~FF  (.D(\u_state_machine/n150 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_state_machine/next_state.WAITING )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/next_state.WAITING~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/next_state.WAITING~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/next_state.WAITING~FF .SR_POLARITY = 1'b1;
    defparam \u_state_machine/next_state.WAITING~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/next_state.WAITING~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/next_state.WAITING~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/next_state.WAITING~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/next_state.WORKING~FF  (.D(\u_state_machine/n150 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_state_machine/next_state.WORKING )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/next_state.WORKING~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/next_state.WORKING~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/next_state.WORKING~FF .SR_POLARITY = 1'b1;
    defparam \u_state_machine/next_state.WORKING~FF .D_POLARITY = 1'b0;
    defparam \u_state_machine/next_state.WORKING~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/next_state.WORKING~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/next_state.WORKING~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/key0_debounced~FF  (.D(\u_state_machine/n5 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_state_machine/key0_debounced )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(28)
    defparam \u_state_machine/key0_debounced~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/key0_debounced~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/key0_debounced~FF .SR_POLARITY = 1'b1;
    defparam \u_state_machine/key0_debounced~FF .D_POLARITY = 1'b0;
    defparam \u_state_machine/key0_debounced~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/key0_debounced~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/key0_debounced~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[1]~FF  (.D(\u_state_machine/n112 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[1]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[1]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[1]~FF .D_POLARITY = 1'b1;
    defparam \led_data[1]~FF .SR_SYNC = 1'b1;
    defparam \led_data[1]~FF .SR_VALUE = 1'b0;
    defparam \led_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[2]~FF  (.D(\u_state_machine/n111 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[2]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[2]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[2]~FF .D_POLARITY = 1'b1;
    defparam \led_data[2]~FF .SR_SYNC = 1'b1;
    defparam \led_data[2]~FF .SR_VALUE = 1'b0;
    defparam \led_data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[3]~FF  (.D(\u_state_machine/n110 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[3]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[3]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[3]~FF .D_POLARITY = 1'b1;
    defparam \led_data[3]~FF .SR_SYNC = 1'b1;
    defparam \led_data[3]~FF .SR_VALUE = 1'b0;
    defparam \led_data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[4]~FF  (.D(\u_state_machine/n109 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[4]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[4]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[4]~FF .D_POLARITY = 1'b1;
    defparam \led_data[4]~FF .SR_SYNC = 1'b1;
    defparam \led_data[4]~FF .SR_VALUE = 1'b0;
    defparam \led_data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[5]~FF  (.D(\u_state_machine/n108 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[5]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[5]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[5]~FF .D_POLARITY = 1'b1;
    defparam \led_data[5]~FF .SR_SYNC = 1'b1;
    defparam \led_data[5]~FF .SR_VALUE = 1'b0;
    defparam \led_data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[6]~FF  (.D(\u_state_machine/n107 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[6]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[6]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[6]~FF .D_POLARITY = 1'b1;
    defparam \led_data[6]~FF .SR_SYNC = 1'b1;
    defparam \led_data[6]~FF .SR_VALUE = 1'b0;
    defparam \led_data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data[7]~FF  (.D(\u_state_machine/n106 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(led_data[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \led_data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \led_data[7]~FF .CE_POLARITY = 1'b1;
    defparam \led_data[7]~FF .SR_POLARITY = 1'b1;
    defparam \led_data[7]~FF .D_POLARITY = 1'b1;
    defparam \led_data[7]~FF .SR_SYNC = 1'b1;
    defparam \led_data[7]~FF .SR_VALUE = 1'b0;
    defparam \led_data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[1]~FF  (.D(\u_state_machine/n98 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[1]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[1]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[1]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[2]~FF  (.D(\u_state_machine/n97 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[2]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[2]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[2]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[3]~FF  (.D(\u_state_machine/n96 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[3]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[3]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[3]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[4]~FF  (.D(\u_state_machine/n95 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[4]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[4]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[4]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[5]~FF  (.D(\u_state_machine/n94 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[5]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[5]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[5]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[6]~FF  (.D(\u_state_machine/n93 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[6]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[6]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[6]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[7]~FF  (.D(\u_state_machine/n92 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[7]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[7]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[7]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[8]~FF  (.D(\u_state_machine/n91 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[8]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[8]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[8]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[9]~FF  (.D(\u_state_machine/n90 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[9]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[9]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[9]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[10]~FF  (.D(\u_state_machine/n89 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[10]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[10]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[10]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[11]~FF  (.D(\u_state_machine/n88 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[11]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[11]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[11]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[12]~FF  (.D(\u_state_machine/n87 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[12]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[12]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[12]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[13]~FF  (.D(\u_state_machine/n86 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[13]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[13]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[13]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[14]~FF  (.D(\u_state_machine/n85 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[14]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[14]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[14]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[15]~FF  (.D(\u_state_machine/n84 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[15]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[15]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[15]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[16]~FF  (.D(\u_state_machine/n83 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[16]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[16]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[16]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[17]~FF  (.D(\u_state_machine/n82 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[17]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[17]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[17]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[18]~FF  (.D(\u_state_machine/n81 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[18]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[18]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[18]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[19]~FF  (.D(\u_state_machine/n80 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[19]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[19]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[19]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[20]~FF  (.D(\u_state_machine/n79 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[20]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[20]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[20]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[20]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[21]~FF  (.D(\u_state_machine/n78 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[21]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[21]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[21]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[21]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[22]~FF  (.D(\u_state_machine/n77 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[22]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[22]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[22]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[22]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[23]~FF  (.D(\u_state_machine/n76 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[23]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[23]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[23]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[23]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[24]~FF  (.D(\u_state_machine/n75 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[24]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[24]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[24]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[24]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[25]~FF  (.D(\u_state_machine/n74 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[25]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[25]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[25]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[25]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_state_machine/counter_10s[26]~FF  (.D(\u_state_machine/n73 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_state_machine/equal_19/n3 ), 
           .Q(\u_state_machine/counter_10s[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\state_machine.v(61)
    defparam \u_state_machine/counter_10s[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[26]~FF .SR_POLARITY = 1'b0;
    defparam \u_state_machine/counter_10s[26]~FF .D_POLARITY = 1'b1;
    defparam \u_state_machine/counter_10s[26]~FF .SR_SYNC = 1'b1;
    defparam \u_state_machine/counter_10s[26]~FF .SR_VALUE = 1'b0;
    defparam \u_state_machine/counter_10s[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__13702 (.I0(\DdrCtrl_ARADDR_0[22] ), .I1(\DdrCtrl_AWADDR_0[22] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13702.LUTMASK = 16'hcaca;
    EFX_FF \w_hdmi_txd0[0]~FF  (.D(\u_rgb2dvi/enc_0/n869 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[0]~FF  (.D(n3464), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_0/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[4]~FF  (.D(\u_rgb2dvi/enc_0/n770 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[8]~FF  (.D(\u_rgb2dvi/enc_0/n806 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[8]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[9]~FF  (.D(\u_rgb2dvi/enc_0/n812 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[1]~FF  (.D(n2836), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_0/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[2]~FF  (.D(n2834), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_0/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[3]~FF  (.D(n2832), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_0/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[4]~FF  (.D(n2831), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_0/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[0]~FF  (.D(\u_rgb2dvi/enc_1/acc[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_lcd_driver/r_lcd_dv ), .Q(\w_hdmi_txd1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[0]~FF  (.D(n3478), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_1/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[4]~FF  (.D(\u_rgb2dvi/enc_1/acc[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_lcd_driver/r_lcd_dv ), .Q(\w_hdmi_txd1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[8]~FF  (.D(n7221), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\w_hdmi_txd1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[8]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[9]~FF  (.D(\u_rgb2dvi/enc_1/q_out[9] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_lcd_driver/r_lcd_dv ), .Q(\w_hdmi_txd1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[1]~FF  (.D(n2786), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_1/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[2]~FF  (.D(n2784), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_1/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[3]~FF  (.D(n2782), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_1/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[4]~FF  (.D(n2781), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_1/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[0]~FF  (.D(\u_rgb2dvi/enc_2/acc[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_lcd_driver/r_lcd_dv ), .Q(\w_hdmi_txd2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[0]~FF  (.D(n3490), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_2/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[4]~FF  (.D(\u_rgb2dvi/enc_2/acc[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_lcd_driver/r_lcd_dv ), .Q(\w_hdmi_txd2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[9]~FF  (.D(\u_rgb2dvi/enc_2/q_out[9] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_lcd_driver/r_lcd_dv ), .Q(\w_hdmi_txd2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[1]~FF  (.D(n2777), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_2/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[2]~FF  (.D(n2775), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_2/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[3]~FF  (.D(n2773), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_2/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[4]~FF  (.D(n2772), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_lcd_driver/r_lcd_dv ), .Q(\u_rgb2dvi/enc_2/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_txc_o[4]~FF  (.D(\r_hdmi_txc_o[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(hdmi_txc_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_txc_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_txc_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_txc_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_txc_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_txc_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_txc_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_txc_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_txc_o[9]~FF  (.D(rc_hdmi_tx), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(\r_hdmi_txc_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_txc_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_txc_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[1]~FF  (.D(n926_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx0_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[2]~FF  (.D(n925_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx0_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[3]~FF  (.D(n924_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx0_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[4]~FF  (.D(n923_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx0_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[6]~FF  (.D(\w_hdmi_txd0[4] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx0_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[7]~FF  (.D(\w_hdmi_txd0[0] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx0_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[8]~FF  (.D(\w_hdmi_txd0[8] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx0_o[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[9]~FF  (.D(\w_hdmi_txd0[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx0_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[1]~FF  (.D(n937_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx1_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[2]~FF  (.D(n936_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx1_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[3]~FF  (.D(n935_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx1_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[4]~FF  (.D(n934_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx1_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[6]~FF  (.D(\w_hdmi_txd1[4] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx1_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[7]~FF  (.D(\w_hdmi_txd1[0] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx1_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[8]~FF  (.D(\w_hdmi_txd1[8] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx1_o[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[9]~FF  (.D(\w_hdmi_txd1[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx1_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[1]~FF  (.D(n948_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx2_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[2]~FF  (.D(n947_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx2_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[3]~FF  (.D(n946_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx2_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[4]~FF  (.D(n945_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \hdmi_tx2_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[6]~FF  (.D(\w_hdmi_txd2[4] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx2_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[7]~FF  (.D(\w_hdmi_txd2[0] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx2_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[9]~FF  (.D(\w_hdmi_txd2[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(700)
    defparam \r_hdmi_tx2_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[1]~FF  (.D(n32_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[2]~FF  (.D(n31_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[3]~FF  (.D(n30_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[4]~FF  (.D(n29_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[5]~FF  (.D(n28_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[6]~FF  (.D(n27_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[7]~FF  (.D(n26_2), .CE(1'b1), .CLK(\Axi0Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(224)
    defparam \PowerOnResetCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \add_82/i4  (.I0(n629), .I1(n654), .CI(1'b0), .O(n405), 
            .CO(n406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i4 .I0_POLARITY = 1'b1;
    defparam \add_82/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i4  (.I0(n405), .I1(n694), .CI(1'b0), .CO(n419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i4 .I0_POLARITY = 1'b1;
    defparam \add_84/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(1'b0), .CI(n12141), .O(n420), .CO(n421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i1  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[0] ), .CI(1'b0), .O(n431), 
            .CO(n432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i1 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i1  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[0] ), .CI(1'b0), .O(n453), 
            .CO(n454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i1 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i1  (.I0(\i2c_config_index[1] ), 
            .I1(\i2c_config_index[0] ), .CI(1'b0), .O(n456), .CO(n457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i1 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i1  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[1] ), .I1(\u_Sensor_Image_XYCrop_0/image_xpos[0] ), 
            .CI(1'b0), .O(n463), .CO(n464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i1 .I0_POLARITY = 1'b1;
    defparam \add_214/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i7  (.I0(n626), .I1(n651), .CI(n1650), .O(n501), 
            .CO(n502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i7 .I0_POLARITY = 1'b1;
    defparam \add_82/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i1  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[1] ), 
            .I1(\u_Sensor_Image_XYCrop_0/image_ypos[0] ), .CI(1'b0), .O(n541), 
            .CO(n542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i1 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i1  (.I0(\u_axi4_ctrl_0/rc_burst[0] ), .I1(DdrCtrl_WREADY_0), 
            .CI(1'b0), .O(n546), .CO(n547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i2  (.I0(\DdrCtrl_ARADDR_0[10] ), .I1(1'b0), 
            .CI(n1197), .O(n631), .CO(n632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i1  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n929), .CO(n930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i2  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n930), .O(n954), .CO(n955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i1  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n958), .CO(n959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] ), .CI(n12142), 
            .O(n961), .CO(n962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i1  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] ), 
            .I1(n5390), .CI(n12143), .CO(n977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/sub_131/add_2/i1  (.I0(\u_axi4_ctrl_0/rfifo_cnt[0] ), 
            .I1(1'b0), .CI(n12144), .O(n978), .CO(n979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(356)
    defparam \u_axi4_ctrl_0/sub_131/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/sub_131/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i1  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n1194), .CO(n1195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i1  (.I0(\DdrCtrl_ARADDR_0[9] ), .I1(\DdrCtrl_ARADDR_0[8] ), 
            .CI(1'b0), .O(n1196), .CO(n1197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i2  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n1195), .O(n1201), .CO(n1202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i1  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n1205), .CO(n1206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] ), .CI(n12145), 
            .O(n1208), .CO(n1209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i1  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] ), 
            .CI(n12146), .CO(n1225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_lcd_driver/add_77/i1  (.I0(\u_lcd_driver/hcnt[1] ), .I1(\u_lcd_driver/hcnt[0] ), 
            .CI(1'b0), .O(n1479), .CO(n1480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i1 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i6  (.I0(n627), .I1(n652), .CI(n1652), .O(n1649), 
            .CO(n1650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i6 .I0_POLARITY = 1'b1;
    defparam \add_82/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i5  (.I0(n628), .I1(n653), .CI(n406), .O(n1651), 
            .CO(n1652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i5 .I0_POLARITY = 1'b1;
    defparam \add_82/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i1  (.I0(\u_lcd_driver/vcnt[1] ), .I1(\u_lcd_driver/vcnt[0] ), 
            .CI(1'b0), .O(n1653), .CO(n1654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i1 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i2  (.I0(\u_lcd_driver/hcnt[1] ), .I1(1'b0), 
            .CI(n12148), .O(n1657), .CO(n1658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i1  (.I0(\u_lcd_driver/vcnt[0] ), .I1(1'b0), 
            .CI(n12149), .O(n1662), .CO(n1663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i1  (.I0(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(1'b0), .O(n1679), 
            .CO(n1680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i1 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i1  (.I0(\u_black_pixel_avg/x_sum[0] ), 
            .I1(\lcd_xpos[0] ), .CI(1'b0), .O(n1714), .CO(n1715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i1 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i1  (.I0(\u_black_pixel_avg/y_sum[0] ), 
            .I1(\lcd_ypos[0] ), .CI(1'b0), .O(n1716), .CO(n1717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i1 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i8  (.I0(\PowerOnResetCnt[7] ), .I1(1'b0), .CI(n1726), 
            .O(n1724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i8 .I0_POLARITY = 1'b1;
    defparam \add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i7  (.I0(\PowerOnResetCnt[6] ), .I1(1'b0), .CI(n1728), 
            .O(n1725), .CO(n1726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i7 .I0_POLARITY = 1'b1;
    defparam \add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i6  (.I0(\PowerOnResetCnt[5] ), .I1(1'b0), .CI(n1730), 
            .O(n1727), .CO(n1728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i6 .I0_POLARITY = 1'b1;
    defparam \add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i5  (.I0(\PowerOnResetCnt[4] ), .I1(1'b0), .CI(n1732), 
            .O(n1729), .CO(n1730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i5 .I0_POLARITY = 1'b1;
    defparam \add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i4  (.I0(\PowerOnResetCnt[3] ), .I1(1'b0), .CI(n1734), 
            .O(n1731), .CO(n1732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i4 .I0_POLARITY = 1'b1;
    defparam \add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i3  (.I0(\PowerOnResetCnt[2] ), .I1(1'b0), .CI(n1736), 
            .O(n1733), .CO(n1734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i3 .I0_POLARITY = 1'b1;
    defparam \add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i2  (.I0(\PowerOnResetCnt[1] ), .I1(1'b0), .CI(n1738), 
            .O(n1735), .CO(n1736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i2 .I0_POLARITY = 1'b1;
    defparam \add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i1  (.I0(\PowerOnResetCnt[0] ), .I1(\reduce_nand_9/n7 ), 
            .CI(1'b0), .O(n1737), .CO(n1738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(223)
    defparam \add_10/i1 .I0_POLARITY = 1'b1;
    defparam \add_10/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_198/i32  (.I0(\u_black_pixel_avg/x_sum[31] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12150), 
            .O(n1812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_198/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_198/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_326/i32  (.I0(n6202), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1815), .O(n1813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_326/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_326/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_326/i31  (.I0(\u_black_pixel_avg/x_sum[30] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12151), 
            .O(n1814), .CO(n1815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_326/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_326/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_452/i32  (.I0(n6206), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1818), .O(n1816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_452/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_452/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_452/i31  (.I0(n6209), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1820), .O(n1817), .CO(n1818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_452/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_452/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_452/i30  (.I0(\u_black_pixel_avg/x_sum[29] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12152), 
            .O(n1819), .CO(n1820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_452/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_452/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_576/i32  (.I0(n6212), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1823), .O(n1821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_576/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_576/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_576/i31  (.I0(n6215), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1825), .O(n1822), .CO(n1823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_576/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_576/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_576/i30  (.I0(n6217), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1827), .O(n1824), .CO(n1825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_576/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_576/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_576/i29  (.I0(\u_black_pixel_avg/x_sum[28] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12153), 
            .O(n1826), .CO(n1827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_576/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_576/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_698/i32  (.I0(n6220), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1830), .O(n1828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_698/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_698/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_698/i31  (.I0(n6223), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1832), .O(n1829), .CO(n1830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_698/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_698/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_698/i30  (.I0(n6225), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1834), .O(n1831), .CO(n1832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_698/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_698/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_698/i29  (.I0(n6227), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1836), .O(n1833), .CO(n1834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_698/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_698/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_698/i28  (.I0(\u_black_pixel_avg/x_sum[27] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12154), 
            .O(n1835), .CO(n1836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_698/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_698/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_818/i32  (.I0(n6230), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1839), .O(n1837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_818/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_818/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_818/i31  (.I0(n6233), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1841), .O(n1838), .CO(n1839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_818/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_818/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_818/i30  (.I0(n6235), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1843), .O(n1840), .CO(n1841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_818/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_818/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_818/i29  (.I0(n6237), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1845), .O(n1842), .CO(n1843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_818/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_818/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_818/i28  (.I0(n6239), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1847), .O(n1844), .CO(n1845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_818/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_818/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_818/i27  (.I0(\u_black_pixel_avg/x_sum[26] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12155), 
            .O(n1846), .CO(n1847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_818/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_818/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_936/i32  (.I0(n6242), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1850), .O(n1848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_936/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_936/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_936/i31  (.I0(n6245), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1852), .O(n1849), .CO(n1850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_936/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_936/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_936/i30  (.I0(n6247), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1854), .O(n1851), .CO(n1852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_936/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_936/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_936/i29  (.I0(n6249), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1856), .O(n1853), .CO(n1854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_936/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_936/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_936/i28  (.I0(n6251), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1858), .O(n1855), .CO(n1856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_936/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_936/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_936/i27  (.I0(n6253), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1860), .O(n1857), .CO(n1858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_936/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_936/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_936/i26  (.I0(\u_black_pixel_avg/x_sum[25] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12156), 
            .O(n1859), .CO(n1860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_936/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_936/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i32  (.I0(n6256), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n1863), .O(n1861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i31  (.I0(n6259), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1865), .O(n1862), .CO(n1863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i30  (.I0(n6261), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1867), .O(n1864), .CO(n1865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i29  (.I0(n6263), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1869), .O(n1866), .CO(n1867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i28  (.I0(n6265), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1871), .O(n1868), .CO(n1869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i27  (.I0(n6267), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1873), .O(n1870), .CO(n1871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i26  (.I0(n6269), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1875), .O(n1872), .CO(n1873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1052/i25  (.I0(\u_black_pixel_avg/x_sum[24] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12157), 
            .O(n1874), .CO(n1875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1052/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1052/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i32  (.I0(n6272), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n1878), .O(n1876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i31  (.I0(n6275), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n1880), .O(n1877), .CO(n1878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i30  (.I0(n6277), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1882), .O(n1879), .CO(n1880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i29  (.I0(n6279), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1884), .O(n1881), .CO(n1882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i28  (.I0(n6281), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1886), .O(n1883), .CO(n1884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i27  (.I0(n6283), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1888), .O(n1885), .CO(n1886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i26  (.I0(n6285), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1890), .O(n1887), .CO(n1888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i25  (.I0(n6287), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1892), .O(n1889), .CO(n1890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1166/i24  (.I0(\u_black_pixel_avg/x_sum[23] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12158), 
            .O(n1891), .CO(n1892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1166/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1166/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i32  (.I0(n6290), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n1895), .O(n1893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i31  (.I0(n6293), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n1897), .O(n1894), .CO(n1895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i30  (.I0(n6295), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n1899), .O(n1896), .CO(n1897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i29  (.I0(n6297), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1901), .O(n1898), .CO(n1899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i28  (.I0(n6299), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1903), .O(n1900), .CO(n1901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i27  (.I0(n6301), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1905), .O(n1902), .CO(n1903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i26  (.I0(n6303), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1907), .O(n1904), .CO(n1905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i25  (.I0(n6305), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1909), .O(n1906), .CO(n1907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i24  (.I0(n6307), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1911), .O(n1908), .CO(n1909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1278/i23  (.I0(\u_black_pixel_avg/x_sum[22] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12159), 
            .O(n1910), .CO(n1911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1278/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1278/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i32  (.I0(n6310), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n1914), .O(n1912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i31  (.I0(n6313), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n1916), .O(n1913), .CO(n1914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i30  (.I0(n6315), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n1918), .O(n1915), .CO(n1916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i29  (.I0(n6317), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n1920), .O(n1917), .CO(n1918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i28  (.I0(n6319), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1922), .O(n1919), .CO(n1920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i27  (.I0(n6321), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1924), .O(n1921), .CO(n1922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i26  (.I0(n6323), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1926), .O(n1923), .CO(n1924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i25  (.I0(n6325), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1928), .O(n1925), .CO(n1926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i24  (.I0(n6327), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1930), .O(n1927), .CO(n1928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i23  (.I0(n6329), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1932), .O(n1929), .CO(n1930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1388/i22  (.I0(\u_black_pixel_avg/x_sum[21] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12160), 
            .O(n1931), .CO(n1932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1388/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1388/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i32  (.I0(n6332), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n1935), .O(n1933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i31  (.I0(n6335), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n1937), .O(n1934), .CO(n1935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i30  (.I0(n6337), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n1939), .O(n1936), .CO(n1937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i29  (.I0(n6339), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n1941), .O(n1938), .CO(n1939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i28  (.I0(n6341), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n1943), .O(n1940), .CO(n1941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i27  (.I0(n6343), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1945), .O(n1942), .CO(n1943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i26  (.I0(n6345), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1947), .O(n1944), .CO(n1945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i25  (.I0(n6347), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1949), .O(n1946), .CO(n1947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i24  (.I0(n6349), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1951), .O(n1948), .CO(n1949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i23  (.I0(n6351), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1953), .O(n1950), .CO(n1951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i22  (.I0(n6353), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1955), .O(n1952), .CO(n1953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1496/i21  (.I0(\u_black_pixel_avg/x_sum[20] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12161), 
            .O(n1954), .CO(n1955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1496/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1496/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i32  (.I0(n6356), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n1958), .O(n1956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i31  (.I0(n6359), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n1960), .O(n1957), .CO(n1958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i30  (.I0(n6361), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n1962), .O(n1959), .CO(n1960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i29  (.I0(n6363), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n1964), .O(n1961), .CO(n1962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i28  (.I0(n6365), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n1966), .O(n1963), .CO(n1964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i27  (.I0(n6367), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n1968), .O(n1965), .CO(n1966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i26  (.I0(n6369), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1970), .O(n1967), .CO(n1968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i25  (.I0(n6371), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1972), .O(n1969), .CO(n1970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i24  (.I0(n6373), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n1974), .O(n1971), .CO(n1972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i23  (.I0(n6375), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n1976), .O(n1973), .CO(n1974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i22  (.I0(n6377), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n1978), .O(n1975), .CO(n1976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i21  (.I0(n6379), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n1980), .O(n1977), .CO(n1978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1602/i20  (.I0(\u_black_pixel_avg/x_sum[19] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12162), 
            .O(n1979), .CO(n1980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1602/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1602/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i32  (.I0(n6382), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n1983), .O(n1981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i31  (.I0(n6385), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n1985), .O(n1982), .CO(n1983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i30  (.I0(n6387), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n1987), .O(n1984), .CO(n1985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i29  (.I0(n6389), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n1989), .O(n1986), .CO(n1987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i28  (.I0(n6391), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n1991), .O(n1988), .CO(n1989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i27  (.I0(n6393), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n1993), .O(n1990), .CO(n1991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i26  (.I0(n6395), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n1995), .O(n1992), .CO(n1993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i25  (.I0(n6397), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n1997), .O(n1994), .CO(n1995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i24  (.I0(n6399), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n1999), .O(n1996), .CO(n1997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i23  (.I0(n6401), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2001), .O(n1998), .CO(n1999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i22  (.I0(n6403), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2003), .O(n2000), .CO(n2001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i21  (.I0(n6405), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2005), .O(n2002), .CO(n2003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i20  (.I0(n6407), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2007), .O(n2004), .CO(n2005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1706/i19  (.I0(\u_black_pixel_avg/x_sum[18] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12163), 
            .O(n2006), .CO(n2007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1706/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1706/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i32  (.I0(n6410), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2010), .O(n2008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i31  (.I0(n6413), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2012), .O(n2009), .CO(n2010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i30  (.I0(n6415), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2014), .O(n2011), .CO(n2012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i29  (.I0(n6417), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2016), .O(n2013), .CO(n2014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i28  (.I0(n6419), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2018), .O(n2015), .CO(n2016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i27  (.I0(n6421), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2020), .O(n2017), .CO(n2018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i26  (.I0(n6423), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2022), .O(n2019), .CO(n2020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i25  (.I0(n6425), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2024), .O(n2021), .CO(n2022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i24  (.I0(n6427), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2026), .O(n2023), .CO(n2024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i23  (.I0(n6429), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2028), .O(n2025), .CO(n2026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i22  (.I0(n6431), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2030), .O(n2027), .CO(n2028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i21  (.I0(n6433), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2032), .O(n2029), .CO(n2030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i20  (.I0(n6435), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2034), .O(n2031), .CO(n2032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i19  (.I0(n6437), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2036), .O(n2033), .CO(n2034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1808/i18  (.I0(\u_black_pixel_avg/x_sum[17] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12164), 
            .O(n2035), .CO(n2036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1808/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1808/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i32  (.I0(n6440), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2039), .O(n2037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i31  (.I0(n6443), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2041), .O(n2038), .CO(n2039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i30  (.I0(n6445), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2043), .O(n2040), .CO(n2041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i29  (.I0(n6447), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2045), .O(n2042), .CO(n2043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i28  (.I0(n6449), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2047), .O(n2044), .CO(n2045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i27  (.I0(n6451), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2049), .O(n2046), .CO(n2047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i26  (.I0(n6453), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2051), .O(n2048), .CO(n2049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i25  (.I0(n6455), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2053), .O(n2050), .CO(n2051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i24  (.I0(n6457), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2055), .O(n2052), .CO(n2053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i23  (.I0(n6459), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2057), .O(n2054), .CO(n2055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i22  (.I0(n6461), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2059), .O(n2056), .CO(n2057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i21  (.I0(n6463), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2061), .O(n2058), .CO(n2059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i20  (.I0(n6465), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2063), .O(n2060), .CO(n2061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i19  (.I0(n6467), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2065), .O(n2062), .CO(n2063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i18  (.I0(n6469), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2067), .O(n2064), .CO(n2065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_1908/i17  (.I0(\u_black_pixel_avg/x_sum[16] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12165), 
            .O(n2066), .CO(n2067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_1908/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_1908/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i32  (.I0(n6472), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n2070), .O(n2068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i31  (.I0(n6475), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2072), .O(n2069), .CO(n2070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i30  (.I0(n6477), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2074), .O(n2071), .CO(n2072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i29  (.I0(n6479), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2076), .O(n2073), .CO(n2074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i28  (.I0(n6481), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2078), .O(n2075), .CO(n2076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i27  (.I0(n6483), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2080), .O(n2077), .CO(n2078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i26  (.I0(n6485), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2082), .O(n2079), .CO(n2080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i25  (.I0(n6487), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2084), .O(n2081), .CO(n2082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i24  (.I0(n6489), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2086), .O(n2083), .CO(n2084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i23  (.I0(n6491), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2088), .O(n2085), .CO(n2086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i22  (.I0(n6493), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2090), .O(n2087), .CO(n2088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i21  (.I0(n6495), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2092), .O(n2089), .CO(n2090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i20  (.I0(n6497), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2094), .O(n2091), .CO(n2092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i19  (.I0(n6499), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2096), .O(n2093), .CO(n2094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i18  (.I0(n6501), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2098), .O(n2095), .CO(n2096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i17  (.I0(n6503), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2100), .O(n2097), .CO(n2098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2006/i16  (.I0(\u_black_pixel_avg/x_sum[15] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12166), 
            .O(n2099), .CO(n2100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2006/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2006/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i30  (.I0(n6506), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2104), .O(n2101), .CO(n2102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i29  (.I0(n6508), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2106), .O(n2103), .CO(n2104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i28  (.I0(n6510), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2108), .O(n2105), .CO(n2106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i27  (.I0(n6512), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2110), .O(n2107), .CO(n2108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i26  (.I0(n6514), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2112), .O(n2109), .CO(n2110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i25  (.I0(n6516), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2114), .O(n2111), .CO(n2112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i24  (.I0(n6518), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2116), .O(n2113), .CO(n2114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i23  (.I0(n6520), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2118), .O(n2115), .CO(n2116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i22  (.I0(n6522), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2120), .O(n2117), .CO(n2118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i21  (.I0(n6524), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2122), .O(n2119), .CO(n2120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i20  (.I0(n6526), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2124), .O(n2121), .CO(n2122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i19  (.I0(n6528), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2126), .O(n2123), .CO(n2124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i18  (.I0(n6530), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2128), .O(n2125), .CO(n2126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i17  (.I0(n6532), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2130), .O(n2127), .CO(n2128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i16  (.I0(n6534), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2132), .O(n2129), .CO(n2130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i15  (.I0(\u_black_pixel_avg/x_sum[14] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12167), 
            .O(n2131), .CO(n2132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i28  (.I0(n6537), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2136), .O(n2133), .CO(n2134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i27  (.I0(n6539), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2138), .O(n2135), .CO(n2136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i26  (.I0(n6541), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2140), .O(n2137), .CO(n2138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i25  (.I0(n6543), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2142), .O(n2139), .CO(n2140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i24  (.I0(n6545), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2144), .O(n2141), .CO(n2142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i23  (.I0(n6547), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2146), .O(n2143), .CO(n2144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i22  (.I0(n6549), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2148), .O(n2145), .CO(n2146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i21  (.I0(n6551), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2150), .O(n2147), .CO(n2148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i20  (.I0(n6553), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2152), .O(n2149), .CO(n2150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i19  (.I0(n6555), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2154), .O(n2151), .CO(n2152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i18  (.I0(n6557), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2156), .O(n2153), .CO(n2154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i17  (.I0(n6559), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2158), .O(n2155), .CO(n2156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i16  (.I0(n6561), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2160), .O(n2157), .CO(n2158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i15  (.I0(n6563), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2162), .O(n2159), .CO(n2160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i14  (.I0(\u_black_pixel_avg/x_sum[13] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12168), 
            .O(n2161), .CO(n2162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i26  (.I0(n6566), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2166), .O(n2163), .CO(n2164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i25  (.I0(n6568), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2168), .O(n2165), .CO(n2166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i24  (.I0(n6570), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2170), .O(n2167), .CO(n2168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i23  (.I0(n6572), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2172), .O(n2169), .CO(n2170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i22  (.I0(n6574), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2174), .O(n2171), .CO(n2172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i21  (.I0(n6576), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2176), .O(n2173), .CO(n2174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i20  (.I0(n6578), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2178), .O(n2175), .CO(n2176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i19  (.I0(n6580), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2180), .O(n2177), .CO(n2178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i18  (.I0(n6582), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2182), .O(n2179), .CO(n2180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i17  (.I0(n6584), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2184), .O(n2181), .CO(n2182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i16  (.I0(n6586), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2186), .O(n2183), .CO(n2184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i15  (.I0(n6588), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2188), .O(n2185), .CO(n2186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i14  (.I0(n6590), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2190), .O(n2187), .CO(n2188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i13  (.I0(\u_black_pixel_avg/x_sum[12] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12169), 
            .O(n2189), .CO(n2190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i24  (.I0(n6593), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2194), .O(n2191), .CO(n2192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i23  (.I0(n6595), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2196), .O(n2193), .CO(n2194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i22  (.I0(n6597), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2198), .O(n2195), .CO(n2196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i21  (.I0(n6599), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2200), .O(n2197), .CO(n2198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i20  (.I0(n6601), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2202), .O(n2199), .CO(n2200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i19  (.I0(n6603), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2204), .O(n2201), .CO(n2202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i18  (.I0(n6605), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2206), .O(n2203), .CO(n2204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i17  (.I0(n6607), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2208), .O(n2205), .CO(n2206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i16  (.I0(n6609), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2210), .O(n2207), .CO(n2208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i15  (.I0(n6611), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2212), .O(n2209), .CO(n2210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i14  (.I0(n6613), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2214), .O(n2211), .CO(n2212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i13  (.I0(n6615), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2216), .O(n2213), .CO(n2214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i12  (.I0(\u_black_pixel_avg/x_sum[11] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12170), 
            .O(n2215), .CO(n2216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i22  (.I0(n6618), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2220), .O(n2217), .CO(n2218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i21  (.I0(n6620), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2222), .O(n2219), .CO(n2220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i20  (.I0(n6622), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2224), .O(n2221), .CO(n2222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i19  (.I0(n6624), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2226), .O(n2223), .CO(n2224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i18  (.I0(n6626), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2228), .O(n2225), .CO(n2226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i17  (.I0(n6628), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2230), .O(n2227), .CO(n2228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i16  (.I0(n6630), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2232), .O(n2229), .CO(n2230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i15  (.I0(n6632), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2234), .O(n2231), .CO(n2232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i14  (.I0(n6634), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2236), .O(n2233), .CO(n2234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i13  (.I0(n6636), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2238), .O(n2235), .CO(n2236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i12  (.I0(n6638), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2240), .O(n2237), .CO(n2238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i11  (.I0(\u_black_pixel_avg/x_sum[10] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12171), 
            .O(n2239), .CO(n2240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i20  (.I0(n6641), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2244), .O(n2241), .CO(n2242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i19  (.I0(n6643), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2246), .O(n2243), .CO(n2244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i18  (.I0(n6645), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2248), .O(n2245), .CO(n2246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i17  (.I0(n6647), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2250), .O(n2247), .CO(n2248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i16  (.I0(n6649), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2252), .O(n2249), .CO(n2250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i15  (.I0(n6651), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2254), .O(n2251), .CO(n2252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i14  (.I0(n6653), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2256), .O(n2253), .CO(n2254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i13  (.I0(n6655), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2258), .O(n2255), .CO(n2256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i12  (.I0(n6657), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2260), .O(n2257), .CO(n2258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i11  (.I0(n6659), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2262), .O(n2259), .CO(n2260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i10  (.I0(\u_black_pixel_avg/x_sum[9] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12172), 
            .O(n2261), .CO(n2262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i18  (.I0(n6662), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2266), .O(n2263), .CO(n2264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i17  (.I0(n6664), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2268), .O(n2265), .CO(n2266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i16  (.I0(n6666), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2270), .O(n2267), .CO(n2268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i15  (.I0(n6668), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2272), .O(n2269), .CO(n2270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i14  (.I0(n6670), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2274), .O(n2271), .CO(n2272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i13  (.I0(n6672), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2276), .O(n2273), .CO(n2274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i12  (.I0(n6674), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2278), .O(n2275), .CO(n2276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i11  (.I0(n6676), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2280), .O(n2277), .CO(n2278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i10  (.I0(n6678), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2282), .O(n2279), .CO(n2280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i9  (.I0(\u_black_pixel_avg/x_sum[8] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12173), 
            .O(n2281), .CO(n2282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i16  (.I0(n6681), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2286), .O(n2283), .CO(n2284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i15  (.I0(n6683), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2288), .O(n2285), .CO(n2286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i14  (.I0(n6685), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2290), .O(n2287), .CO(n2288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i13  (.I0(n6687), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2292), .O(n2289), .CO(n2290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i12  (.I0(n6689), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2294), .O(n2291), .CO(n2292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i11  (.I0(n6691), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2296), .O(n2293), .CO(n2294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i10  (.I0(n6693), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2298), .O(n2295), .CO(n2296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i9  (.I0(n6695), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2300), .O(n2297), .CO(n2298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i8  (.I0(\u_black_pixel_avg/x_sum[7] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12174), 
            .O(n2299), .CO(n2300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_198/i32  (.I0(\u_black_pixel_avg/y_sum[31] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12181), 
            .O(n2367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_198/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_198/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_326/i32  (.I0(n6759), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2370), .O(n2368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_326/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_326/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_326/i31  (.I0(\u_black_pixel_avg/y_sum[30] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12182), 
            .O(n2369), .CO(n2370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_326/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_326/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_452/i32  (.I0(n6762), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2373), .O(n2371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_452/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_452/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_452/i31  (.I0(n6764), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2375), .O(n2372), .CO(n2373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_452/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_452/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_452/i30  (.I0(\u_black_pixel_avg/y_sum[29] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12183), 
            .O(n2374), .CO(n2375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_452/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_452/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_576/i32  (.I0(n6767), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2378), .O(n2376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_576/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_576/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_576/i31  (.I0(n6769), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2380), .O(n2377), .CO(n2378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_576/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_576/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_576/i30  (.I0(n6771), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2382), .O(n2379), .CO(n2380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_576/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_576/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_576/i29  (.I0(\u_black_pixel_avg/y_sum[28] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12184), 
            .O(n2381), .CO(n2382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_576/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_576/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_698/i32  (.I0(n6774), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2385), .O(n2383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_698/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_698/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_698/i31  (.I0(n6776), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2387), .O(n2384), .CO(n2385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_698/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_698/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_698/i30  (.I0(n6778), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2389), .O(n2386), .CO(n2387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_698/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_698/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_698/i29  (.I0(n6780), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2391), .O(n2388), .CO(n2389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_698/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_698/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_698/i28  (.I0(\u_black_pixel_avg/y_sum[27] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12185), 
            .O(n2390), .CO(n2391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_698/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_698/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_818/i32  (.I0(n6783), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2394), .O(n2392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_818/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_818/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_818/i31  (.I0(n6785), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2396), .O(n2393), .CO(n2394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_818/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_818/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_818/i30  (.I0(n6787), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2398), .O(n2395), .CO(n2396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_818/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_818/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_818/i29  (.I0(n6789), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2400), .O(n2397), .CO(n2398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_818/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_818/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_818/i28  (.I0(n6791), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2402), .O(n2399), .CO(n2400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_818/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_818/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_818/i27  (.I0(\u_black_pixel_avg/y_sum[26] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12186), 
            .O(n2401), .CO(n2402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_818/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_818/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_936/i32  (.I0(n6794), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2405), .O(n2403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_936/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_936/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_936/i31  (.I0(n6796), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2407), .O(n2404), .CO(n2405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_936/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_936/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_936/i30  (.I0(n6798), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2409), .O(n2406), .CO(n2407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_936/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_936/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_936/i29  (.I0(n6800), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2411), .O(n2408), .CO(n2409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_936/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_936/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_936/i28  (.I0(n6802), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2413), .O(n2410), .CO(n2411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_936/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_936/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_936/i27  (.I0(n6804), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2415), .O(n2412), .CO(n2413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_936/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_936/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_936/i26  (.I0(\u_black_pixel_avg/y_sum[25] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12187), 
            .O(n2414), .CO(n2415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_936/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_936/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i32  (.I0(n6807), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2418), .O(n2416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i31  (.I0(n6809), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2420), .O(n2417), .CO(n2418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i30  (.I0(n6811), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2422), .O(n2419), .CO(n2420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i29  (.I0(n6813), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2424), .O(n2421), .CO(n2422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i28  (.I0(n6815), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2426), .O(n2423), .CO(n2424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i27  (.I0(n6817), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2428), .O(n2425), .CO(n2426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i26  (.I0(n6819), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2430), .O(n2427), .CO(n2428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1052/i25  (.I0(\u_black_pixel_avg/y_sum[24] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12188), 
            .O(n2429), .CO(n2430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1052/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1052/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i32  (.I0(n6822), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2433), .O(n2431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i31  (.I0(n6824), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2435), .O(n2432), .CO(n2433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i30  (.I0(n6826), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2437), .O(n2434), .CO(n2435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i29  (.I0(n6828), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2439), .O(n2436), .CO(n2437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i28  (.I0(n6830), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2441), .O(n2438), .CO(n2439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i27  (.I0(n6832), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2443), .O(n2440), .CO(n2441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i26  (.I0(n6834), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2445), .O(n2442), .CO(n2443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i25  (.I0(n6836), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2447), .O(n2444), .CO(n2445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1166/i24  (.I0(\u_black_pixel_avg/y_sum[23] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12189), 
            .O(n2446), .CO(n2447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1166/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1166/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i32  (.I0(n6839), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2450), .O(n2448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i31  (.I0(n6841), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2452), .O(n2449), .CO(n2450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i30  (.I0(n6843), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2454), .O(n2451), .CO(n2452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i29  (.I0(n6845), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2456), .O(n2453), .CO(n2454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i28  (.I0(n6847), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2458), .O(n2455), .CO(n2456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i27  (.I0(n6849), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2460), .O(n2457), .CO(n2458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i26  (.I0(n6851), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2462), .O(n2459), .CO(n2460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i25  (.I0(n6853), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2464), .O(n2461), .CO(n2462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i24  (.I0(n6855), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2466), .O(n2463), .CO(n2464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1278/i23  (.I0(\u_black_pixel_avg/y_sum[22] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12190), 
            .O(n2465), .CO(n2466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1278/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1278/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i32  (.I0(n6858), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2469), .O(n2467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i31  (.I0(n6860), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2471), .O(n2468), .CO(n2469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i30  (.I0(n6862), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2473), .O(n2470), .CO(n2471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i29  (.I0(n6864), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2475), .O(n2472), .CO(n2473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i28  (.I0(n6866), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2477), .O(n2474), .CO(n2475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i27  (.I0(n6868), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2479), .O(n2476), .CO(n2477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i26  (.I0(n6870), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2481), .O(n2478), .CO(n2479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i25  (.I0(n6872), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2483), .O(n2480), .CO(n2481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i24  (.I0(n6874), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2485), .O(n2482), .CO(n2483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i23  (.I0(n6876), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2487), .O(n2484), .CO(n2485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1388/i22  (.I0(\u_black_pixel_avg/y_sum[21] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12191), 
            .O(n2486), .CO(n2487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1388/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1388/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i32  (.I0(n6879), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2490), .O(n2488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i31  (.I0(n6881), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2492), .O(n2489), .CO(n2490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i30  (.I0(n6883), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2494), .O(n2491), .CO(n2492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i29  (.I0(n6885), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2496), .O(n2493), .CO(n2494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i28  (.I0(n6887), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2498), .O(n2495), .CO(n2496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i27  (.I0(n6889), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2500), .O(n2497), .CO(n2498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i26  (.I0(n6891), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2502), .O(n2499), .CO(n2500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i25  (.I0(n6893), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2504), .O(n2501), .CO(n2502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i24  (.I0(n6895), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2506), .O(n2503), .CO(n2504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i23  (.I0(n6897), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2508), .O(n2505), .CO(n2506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i22  (.I0(n6899), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2510), .O(n2507), .CO(n2508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1496/i21  (.I0(\u_black_pixel_avg/y_sum[20] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12192), 
            .O(n2509), .CO(n2510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1496/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1496/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i32  (.I0(n6902), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2513), .O(n2511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i31  (.I0(n6904), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2515), .O(n2512), .CO(n2513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i30  (.I0(n6906), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2517), .O(n2514), .CO(n2515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i29  (.I0(n6908), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2519), .O(n2516), .CO(n2517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i28  (.I0(n6910), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2521), .O(n2518), .CO(n2519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i27  (.I0(n6912), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2523), .O(n2520), .CO(n2521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i26  (.I0(n6914), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2525), .O(n2522), .CO(n2523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i25  (.I0(n6916), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2527), .O(n2524), .CO(n2525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i24  (.I0(n6918), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2529), .O(n2526), .CO(n2527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i23  (.I0(n6920), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2531), .O(n2528), .CO(n2529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i22  (.I0(n6922), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2533), .O(n2530), .CO(n2531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i21  (.I0(n6924), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2535), .O(n2532), .CO(n2533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1602/i20  (.I0(\u_black_pixel_avg/y_sum[19] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12193), 
            .O(n2534), .CO(n2535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1602/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1602/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i32  (.I0(n6927), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2538), .O(n2536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i31  (.I0(n6929), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2540), .O(n2537), .CO(n2538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i30  (.I0(n6931), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2542), .O(n2539), .CO(n2540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i29  (.I0(n6933), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2544), .O(n2541), .CO(n2542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i28  (.I0(n6935), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2546), .O(n2543), .CO(n2544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i27  (.I0(n6937), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2548), .O(n2545), .CO(n2546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i26  (.I0(n6939), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2550), .O(n2547), .CO(n2548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i25  (.I0(n6941), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2552), .O(n2549), .CO(n2550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i24  (.I0(n6943), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2554), .O(n2551), .CO(n2552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i23  (.I0(n6945), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2556), .O(n2553), .CO(n2554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i22  (.I0(n6947), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2558), .O(n2555), .CO(n2556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i21  (.I0(n6949), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2560), .O(n2557), .CO(n2558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i20  (.I0(n6951), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2562), .O(n2559), .CO(n2560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1706/i19  (.I0(\u_black_pixel_avg/y_sum[18] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12194), 
            .O(n2561), .CO(n2562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1706/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1706/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i32  (.I0(n6954), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2565), .O(n2563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i31  (.I0(n6956), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2567), .O(n2564), .CO(n2565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i30  (.I0(n6958), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2569), .O(n2566), .CO(n2567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i29  (.I0(n6960), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2571), .O(n2568), .CO(n2569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i28  (.I0(n6962), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2573), .O(n2570), .CO(n2571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i27  (.I0(n6964), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2575), .O(n2572), .CO(n2573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i26  (.I0(n6966), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2577), .O(n2574), .CO(n2575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i25  (.I0(n6968), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2579), .O(n2576), .CO(n2577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i24  (.I0(n6970), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2581), .O(n2578), .CO(n2579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i23  (.I0(n6972), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2583), .O(n2580), .CO(n2581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i22  (.I0(n6974), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2585), .O(n2582), .CO(n2583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i21  (.I0(n6976), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2587), .O(n2584), .CO(n2585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i20  (.I0(n6978), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2589), .O(n2586), .CO(n2587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i19  (.I0(n6980), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2591), .O(n2588), .CO(n2589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1808/i18  (.I0(\u_black_pixel_avg/y_sum[17] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12195), 
            .O(n2590), .CO(n2591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1808/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1808/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i32  (.I0(n6983), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2594), .O(n2592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i31  (.I0(n6985), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2596), .O(n2593), .CO(n2594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i30  (.I0(n6987), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2598), .O(n2595), .CO(n2596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i29  (.I0(n6989), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2600), .O(n2597), .CO(n2598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i28  (.I0(n6991), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2602), .O(n2599), .CO(n2600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i27  (.I0(n6993), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2604), .O(n2601), .CO(n2602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i26  (.I0(n6995), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2606), .O(n2603), .CO(n2604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i25  (.I0(n6997), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2608), .O(n2605), .CO(n2606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i24  (.I0(n6999), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2610), .O(n2607), .CO(n2608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i23  (.I0(n7001), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2612), .O(n2609), .CO(n2610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i22  (.I0(n7003), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2614), .O(n2611), .CO(n2612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i21  (.I0(n7005), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2616), .O(n2613), .CO(n2614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i20  (.I0(n7007), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2618), .O(n2615), .CO(n2616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i19  (.I0(n7009), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2620), .O(n2617), .CO(n2618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i18  (.I0(n7011), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2622), .O(n2619), .CO(n2620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_1908/i17  (.I0(\u_black_pixel_avg/y_sum[16] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12196), 
            .O(n2621), .CO(n2622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_1908/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_1908/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i32  (.I0(n7014), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n2625), .O(n2623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i31  (.I0(n7016), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2627), .O(n2624), .CO(n2625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i30  (.I0(n7018), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2629), .O(n2626), .CO(n2627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i29  (.I0(n7020), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2631), .O(n2628), .CO(n2629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i28  (.I0(n7022), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2633), .O(n2630), .CO(n2631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i27  (.I0(n7024), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2635), .O(n2632), .CO(n2633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i26  (.I0(n7026), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2637), .O(n2634), .CO(n2635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i25  (.I0(n7028), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2639), .O(n2636), .CO(n2637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i24  (.I0(n7030), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2641), .O(n2638), .CO(n2639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i23  (.I0(n7032), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2643), .O(n2640), .CO(n2641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i22  (.I0(n7034), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2645), .O(n2642), .CO(n2643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i21  (.I0(n7036), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2647), .O(n2644), .CO(n2645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i20  (.I0(n7038), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2649), .O(n2646), .CO(n2647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i19  (.I0(n7040), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2651), .O(n2648), .CO(n2649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i18  (.I0(n7042), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2653), .O(n2650), .CO(n2651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i17  (.I0(n7044), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2655), .O(n2652), .CO(n2653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2006/i16  (.I0(\u_black_pixel_avg/y_sum[15] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12197), 
            .O(n2654), .CO(n2655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2006/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2006/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i30  (.I0(n7047), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2659), .O(n2656), .CO(n2657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i29  (.I0(n7049), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2661), .O(n2658), .CO(n2659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i28  (.I0(n7051), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2663), .O(n2660), .CO(n2661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i27  (.I0(n7053), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2665), .O(n2662), .CO(n2663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i26  (.I0(n7055), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2667), .O(n2664), .CO(n2665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i25  (.I0(n7057), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2669), .O(n2666), .CO(n2667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i24  (.I0(n7059), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2671), .O(n2668), .CO(n2669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i23  (.I0(n7061), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2673), .O(n2670), .CO(n2671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i22  (.I0(n7063), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2675), .O(n2672), .CO(n2673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i21  (.I0(n7065), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2677), .O(n2674), .CO(n2675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i20  (.I0(n7067), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2679), .O(n2676), .CO(n2677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i19  (.I0(n7069), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2681), .O(n2678), .CO(n2679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i18  (.I0(n7071), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2683), .O(n2680), .CO(n2681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i17  (.I0(n7073), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2685), .O(n2682), .CO(n2683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i16  (.I0(n7075), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2687), .O(n2684), .CO(n2685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i15  (.I0(\u_black_pixel_avg/y_sum[14] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12198), 
            .O(n2686), .CO(n2687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i28  (.I0(n7078), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2691), .O(n2688), .CO(n2689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i27  (.I0(n7080), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2693), .O(n2690), .CO(n2691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i26  (.I0(n7082), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2695), .O(n2692), .CO(n2693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i25  (.I0(n7084), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2697), .O(n2694), .CO(n2695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i24  (.I0(n7086), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2699), .O(n2696), .CO(n2697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i23  (.I0(n7088), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2701), .O(n2698), .CO(n2699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i22  (.I0(n7090), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2703), .O(n2700), .CO(n2701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i21  (.I0(n7092), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2705), .O(n2702), .CO(n2703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i20  (.I0(n7094), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2707), .O(n2704), .CO(n2705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i19  (.I0(n7096), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2709), .O(n2706), .CO(n2707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i18  (.I0(n7098), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2711), .O(n2708), .CO(n2709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i17  (.I0(n7100), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2713), .O(n2710), .CO(n2711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i16  (.I0(n7102), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2715), .O(n2712), .CO(n2713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i15  (.I0(n7104), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2717), .O(n2714), .CO(n2715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i14  (.I0(\u_black_pixel_avg/y_sum[13] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12199), 
            .O(n2716), .CO(n2717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i26  (.I0(n7107), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2721), .O(n2718), .CO(n2719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i25  (.I0(n7109), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2723), .O(n2720), .CO(n2721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i24  (.I0(n7111), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2725), .O(n2722), .CO(n2723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i23  (.I0(n7113), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2727), .O(n2724), .CO(n2725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i22  (.I0(n7115), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2729), .O(n2726), .CO(n2727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i21  (.I0(n7117), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2731), .O(n2728), .CO(n2729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i20  (.I0(n7119), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2733), .O(n2730), .CO(n2731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i19  (.I0(n7121), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2735), .O(n2732), .CO(n2733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i18  (.I0(n7123), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2737), .O(n2734), .CO(n2735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i17  (.I0(n7125), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2739), .O(n2736), .CO(n2737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i16  (.I0(n7127), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2741), .O(n2738), .CO(n2739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i15  (.I0(n7129), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2743), .O(n2740), .CO(n2741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i14  (.I0(n7131), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2745), .O(n2742), .CO(n2743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i13  (.I0(\u_black_pixel_avg/y_sum[12] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12200), 
            .O(n2744), .CO(n2745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i24  (.I0(n7134), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2749), .O(n2746), .CO(n2747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i23  (.I0(n7136), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2751), .O(n2748), .CO(n2749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i22  (.I0(n7138), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2753), .O(n2750), .CO(n2751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i21  (.I0(n7140), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2755), .O(n2752), .CO(n2753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i20  (.I0(n7142), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2757), .O(n2754), .CO(n2755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i19  (.I0(n7144), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2759), .O(n2756), .CO(n2757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i18  (.I0(n7146), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2761), .O(n2758), .CO(n2759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i17  (.I0(n7148), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2763), .O(n2760), .CO(n2761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i16  (.I0(n7150), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2765), .O(n2762), .CO(n2763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i15  (.I0(n7152), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2767), .O(n2764), .CO(n2765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i14  (.I0(n7154), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2769), .O(n2766), .CO(n2767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i13  (.I0(n7156), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2771), .O(n2768), .CO(n2769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i12  (.I0(\u_black_pixel_avg/y_sum[11] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12201), 
            .O(n2770), .CO(n2771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i5  (.I0(\u_rgb2dvi/enc_2/acc[4] ), .I1(n7160), 
            .CI(n2774), .O(n2772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i4  (.I0(\u_rgb2dvi/enc_2/acc[3] ), .I1(n7163), 
            .CI(n2776), .O(n2773), .CO(n2774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i3  (.I0(\u_rgb2dvi/enc_2/acc[2] ), .I1(n7166), 
            .CI(n2778), .O(n2775), .CO(n2776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i2  (.I0(\u_rgb2dvi/enc_2/acc[1] ), .I1(n7169), 
            .CI(n3491), .O(n2777), .CO(n2778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_75/i4  (.I0(n2818), .I1(1'b0), .CI(n3351), 
            .O(n2779), .CO(n2780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_2/add_75/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_75/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i5  (.I0(\u_rgb2dvi/enc_1/acc[4] ), .I1(n7174), 
            .CI(n2783), .O(n2781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i4  (.I0(\u_rgb2dvi/enc_1/acc[3] ), .I1(n7177), 
            .CI(n2785), .O(n2782), .CO(n2783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i3  (.I0(\u_rgb2dvi/enc_1/acc[2] ), .I1(n7180), 
            .CI(n2787), .O(n2784), .CO(n2785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i2  (.I0(\u_rgb2dvi/enc_1/acc[1] ), .I1(n7183), 
            .CI(n3479), .O(n2786), .CO(n2787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i22  (.I0(n7185), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2791), .O(n2788), .CO(n2789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i21  (.I0(n7187), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2793), .O(n2790), .CO(n2791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i20  (.I0(n7189), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2795), .O(n2792), .CO(n2793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i19  (.I0(n7191), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2797), .O(n2794), .CO(n2795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i18  (.I0(n7193), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2799), .O(n2796), .CO(n2797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i17  (.I0(n7195), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2801), .O(n2798), .CO(n2799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i16  (.I0(n7197), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2803), .O(n2800), .CO(n2801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i15  (.I0(n7199), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2805), .O(n2802), .CO(n2803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i14  (.I0(n7201), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2807), .O(n2804), .CO(n2805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i13  (.I0(n7203), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2809), .O(n2806), .CO(n2807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i12  (.I0(n7205), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2811), .O(n2808), .CO(n2809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i11  (.I0(\u_black_pixel_avg/y_sum[10] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12202), 
            .O(n2810), .CO(n2811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i5  (.I0(n2824), .I1(1'b1), .CI(n2814), 
            .O(n2812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i4  (.I0(n2825), .I1(1'b1), .CI(n2816), 
            .O(n2813), .CO(n2814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i3  (.I0(n2827), .I1(1'b1), .CI(n3469), 
            .O(n2815), .CO(n2816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i5  (.I0(1'b0), .I1(1'b1), .CI(n2819), 
            .O(n2817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i4  (.I0(n7221), .I1(n7221), .CI(n2821), 
            .O(n2818), .CO(n2819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i4 .I0_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i3  (.I0(1'b0), .I1(1'b1), .CI(n2823), 
            .O(n2820), .CO(n2821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i2  (.I0(1'b0), .I1(1'b1), .CI(n12216), 
            .O(n2822), .CO(n2823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i5  (.I0(1'b0), .I1(1'b1), .CI(n2826), 
            .O(n2824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i4  (.I0(n7221), .I1(n7221), .CI(n2828), 
            .O(n2825), .CO(n2826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i3  (.I0(1'b0), .I1(1'b1), .CI(n2830), 
            .O(n2827), .CO(n2828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i2  (.I0(1'b0), .I1(1'b1), .CI(n12215), 
            .O(n2829), .CO(n2830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i5  (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(n7226), 
            .CI(n2833), .O(n2831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i4  (.I0(\u_rgb2dvi/enc_0/acc[3] ), .I1(n7229), 
            .CI(n2835), .O(n2832), .CO(n2833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i3  (.I0(\u_rgb2dvi/enc_0/acc[2] ), .I1(n7232), 
            .CI(n2837), .O(n2834), .CO(n2835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i2  (.I0(\u_rgb2dvi/enc_0/acc[1] ), .I1(n7235), 
            .CI(n3465), .O(n2836), .CO(n2837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i5  (.I0(n2817), .I1(1'b0), .CI(n2780), 
            .O(n2838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i20  (.I0(n7245), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2845), .O(n2842), .CO(n2843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i19  (.I0(n7247), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2847), .O(n2844), .CO(n2845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i18  (.I0(n7249), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2849), .O(n2846), .CO(n2847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i17  (.I0(n7251), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2851), .O(n2848), .CO(n2849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i16  (.I0(n7253), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2853), .O(n2850), .CO(n2851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i15  (.I0(n7255), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2855), .O(n2852), .CO(n2853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i14  (.I0(n7257), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2857), .O(n2854), .CO(n2855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i13  (.I0(n7259), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2859), .O(n2856), .CO(n2857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i12  (.I0(n7261), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2861), .O(n2858), .CO(n2859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i11  (.I0(n7263), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2863), .O(n2860), .CO(n2861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i10  (.I0(\u_black_pixel_avg/y_sum[9] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12203), 
            .O(n2862), .CO(n2863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i18  (.I0(n7334), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2922), .O(n2919), .CO(n2920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i17  (.I0(n7336), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2924), .O(n2921), .CO(n2922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i16  (.I0(n7338), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2926), .O(n2923), .CO(n2924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i15  (.I0(n7340), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2928), .O(n2925), .CO(n2926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i14  (.I0(n7342), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n2930), .O(n2927), .CO(n2928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i13  (.I0(n7344), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n2932), .O(n2929), .CO(n2930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i12  (.I0(n7346), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n2934), .O(n2931), .CO(n2932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i11  (.I0(n7348), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n2936), .O(n2933), .CO(n2934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i10  (.I0(n7350), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n2938), .O(n2935), .CO(n2936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i9  (.I0(\u_black_pixel_avg/y_sum[8] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12204), 
            .O(n2937), .CO(n2938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i16  (.I0(n7407), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n2995), .O(n2992), .CO(n2993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i15  (.I0(n7409), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n2997), .O(n2994), .CO(n2995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i14  (.I0(n7411), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n2999), .O(n2996), .CO(n2997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i13  (.I0(n7413), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n3001), .O(n2998), .CO(n2999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i12  (.I0(n7415), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n3003), .O(n3000), .CO(n3001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i11  (.I0(n7417), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n3005), .O(n3002), .CO(n3003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i10  (.I0(n7419), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n3007), .O(n3004), .CO(n3005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i9  (.I0(n7421), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n3009), .O(n3006), .CO(n3007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i8  (.I0(\u_black_pixel_avg/y_sum[7] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12205), 
            .O(n3008), .CO(n3009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i32  (.I0(n7466), .I1(\u_black_pixel_avg/black_pixel_count[27] ), 
            .CI(n3054), .O(n3052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i31  (.I0(n7468), .I1(\u_black_pixel_avg/black_pixel_count[26] ), 
            .CI(n3056), .O(n3053), .CO(n3054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i30  (.I0(n7470), .I1(\u_black_pixel_avg/black_pixel_count[25] ), 
            .CI(n3058), .O(n3055), .CO(n3056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i29  (.I0(n7472), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .CI(n3060), .O(n3057), .CO(n3058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i28  (.I0(n7474), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .CI(n3078), .O(n3059), .CO(n3060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i14  (.I0(n7476), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n3064), .O(n3061), .CO(n3062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i13  (.I0(n7478), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n3066), .O(n3063), .CO(n3064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i12  (.I0(n7480), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n3068), .O(n3065), .CO(n3066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i11  (.I0(n7482), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n3070), .O(n3067), .CO(n3068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i10  (.I0(n7484), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n3072), .O(n3069), .CO(n3070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i9  (.I0(n7486), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n3074), .O(n3071), .CO(n3072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i8  (.I0(n7488), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n3076), .O(n3073), .CO(n3074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i7  (.I0(\u_black_pixel_avg/y_sum[6] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12206), 
            .O(n3075), .CO(n3076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i7 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i27  (.I0(n7491), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3080), .O(n3077), .CO(n3078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i26  (.I0(n7493), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3082), .O(n3079), .CO(n3080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i25  (.I0(n7495), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3084), .O(n3081), .CO(n3082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i24  (.I0(n7497), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3086), .O(n3083), .CO(n3084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i23  (.I0(n7499), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3088), .O(n3085), .CO(n3086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i22  (.I0(n7501), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3090), .O(n3087), .CO(n3088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i21  (.I0(n7503), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3092), .O(n3089), .CO(n3090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i20  (.I0(n7505), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3094), .O(n3091), .CO(n3092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i19  (.I0(n7507), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3096), .O(n3093), .CO(n3094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i18  (.I0(n7509), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3098), .O(n3095), .CO(n3096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i17  (.I0(n7511), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3100), .O(n3097), .CO(n3098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i16  (.I0(n7513), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n3102), .O(n3099), .CO(n3100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i15  (.I0(n7515), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n3104), .O(n3101), .CO(n3102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i14  (.I0(n7517), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n3106), .O(n3103), .CO(n3104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i13  (.I0(n7519), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n3108), .O(n3105), .CO(n3106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i12  (.I0(n7521), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n3110), .O(n3107), .CO(n3108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i11  (.I0(n7523), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n3188), .O(n3109), .CO(n3110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i32  (.I0(n7525), .I1(\u_black_pixel_avg/black_pixel_count[26] ), 
            .CI(n3113), .O(n3111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i31  (.I0(n7527), .I1(\u_black_pixel_avg/black_pixel_count[25] ), 
            .CI(n3115), .O(n3112), .CO(n3113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i30  (.I0(n7529), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .CI(n3117), .O(n3114), .CO(n3115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i29  (.I0(n7531), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .CI(n3119), .O(n3116), .CO(n3117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i28  (.I0(n7533), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3121), .O(n3118), .CO(n3119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i27  (.I0(n7535), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3123), .O(n3120), .CO(n3121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i26  (.I0(n7537), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3125), .O(n3122), .CO(n3123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i25  (.I0(n7539), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3141), .O(n3124), .CO(n3125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i12  (.I0(n7541), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .CI(n3129), .O(n3126), .CO(n3127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i11  (.I0(n7543), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n3131), .O(n3128), .CO(n3129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i10  (.I0(n7545), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n3133), .O(n3130), .CO(n3131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i9  (.I0(n7547), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n3135), .O(n3132), .CO(n3133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i8  (.I0(n7549), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n3137), .O(n3134), .CO(n3135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i7  (.I0(n7551), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n3139), .O(n3136), .CO(n3137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i7 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i6  (.I0(\u_black_pixel_avg/y_sum[5] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12207), 
            .O(n3138), .CO(n3139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i6 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i24  (.I0(n7554), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3143), .O(n3140), .CO(n3141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i23  (.I0(n7556), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3145), .O(n3142), .CO(n3143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i22  (.I0(n7558), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3147), .O(n3144), .CO(n3145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i21  (.I0(n7560), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3149), .O(n3146), .CO(n3147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i20  (.I0(n7562), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3151), .O(n3148), .CO(n3149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i19  (.I0(n7564), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3153), .O(n3150), .CO(n3151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i18  (.I0(n7566), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3155), .O(n3152), .CO(n3153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i17  (.I0(n7568), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n3157), .O(n3154), .CO(n3155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i16  (.I0(n7570), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n3159), .O(n3156), .CO(n3157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i15  (.I0(n7572), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n3161), .O(n3158), .CO(n3159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i14  (.I0(n7574), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n3163), .O(n3160), .CO(n3161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2876/i13  (.I0(n7576), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .CI(n3127), .O(n3162), .CO(n3163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2876/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2876/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i32  (.I0(n7578), .I1(\u_black_pixel_avg/black_pixel_count[25] ), 
            .CI(n3166), .O(n3164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i31  (.I0(n7580), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .CI(n3168), .O(n3165), .CO(n3166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i30  (.I0(n7582), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .CI(n3170), .O(n3167), .CO(n3168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i29  (.I0(n7584), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3172), .O(n3169), .CO(n3170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i28  (.I0(n7586), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3174), .O(n3171), .CO(n3172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i27  (.I0(n7588), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3176), .O(n3173), .CO(n3174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i26  (.I0(n7590), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3178), .O(n3175), .CO(n3176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i25  (.I0(n7592), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3180), .O(n3177), .CO(n3178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i24  (.I0(n7594), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3182), .O(n3179), .CO(n3180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i23  (.I0(n7596), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3184), .O(n3181), .CO(n3182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i22  (.I0(n7598), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3186), .O(n3183), .CO(n3184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i21  (.I0(n7600), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3200), .O(n3185), .CO(n3186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i10  (.I0(n7602), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .CI(n3190), .O(n3187), .CO(n3188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i9  (.I0(n7604), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .CI(n3192), .O(n3189), .CO(n3190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i8  (.I0(n7606), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .CI(n3194), .O(n3191), .CO(n3192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i7  (.I0(n7608), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .CI(n3196), .O(n3193), .CO(n3194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i7 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i6  (.I0(n7610), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .CI(n3198), .O(n3195), .CO(n3196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i6 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2952/i5  (.I0(\u_black_pixel_avg/y_sum[4] ), 
            .I1(\u_black_pixel_avg/black_pixel_count[0] ), .CI(n12208), 
            .O(n3197), .CO(n3198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2952/i5 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2952/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i20  (.I0(n7613), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3202), .O(n3199), .CO(n3200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i19  (.I0(n7615), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3204), .O(n3201), .CO(n3202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i18  (.I0(n7617), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n3206), .O(n3203), .CO(n3204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i17  (.I0(n7619), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n3208), .O(n3205), .CO(n3206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i16  (.I0(n7621), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n3210), .O(n3207), .CO(n3208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2798/i15  (.I0(n7623), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .CI(n3062), .O(n3209), .CO(n3210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2798/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2798/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i32  (.I0(n7625), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .CI(n3213), .O(n3211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i31  (.I0(n7627), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .CI(n3215), .O(n3212), .CO(n3213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i30  (.I0(n7629), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3217), .O(n3214), .CO(n3215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i29  (.I0(n7631), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3219), .O(n3216), .CO(n3217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i28  (.I0(n7633), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3221), .O(n3218), .CO(n3219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i27  (.I0(n7635), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3223), .O(n3220), .CO(n3221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i26  (.I0(n7637), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3225), .O(n3222), .CO(n3223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i25  (.I0(n7639), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3227), .O(n3224), .CO(n3225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i24  (.I0(n7641), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3229), .O(n3226), .CO(n3227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i23  (.I0(n7643), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3231), .O(n3228), .CO(n3229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i22  (.I0(n7645), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3233), .O(n3230), .CO(n3231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i21  (.I0(n7647), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3235), .O(n3232), .CO(n3233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i20  (.I0(n7649), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3237), .O(n3234), .CO(n3235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i19  (.I0(n7651), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n3239), .O(n3236), .CO(n3237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i18  (.I0(n7653), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n3241), .O(n3238), .CO(n3239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2718/i17  (.I0(n7655), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2993), .O(n3240), .CO(n3241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2718/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2718/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i32  (.I0(n7666), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .CI(n3254), .O(n3252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i31  (.I0(n7668), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3256), .O(n3253), .CO(n3254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i30  (.I0(n7670), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3258), .O(n3255), .CO(n3256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i29  (.I0(n7672), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3260), .O(n3257), .CO(n3258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i28  (.I0(n7674), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3262), .O(n3259), .CO(n3260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i27  (.I0(n7676), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3264), .O(n3261), .CO(n3262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i26  (.I0(n7678), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3266), .O(n3263), .CO(n3264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i25  (.I0(n7680), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3268), .O(n3265), .CO(n3266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i24  (.I0(n7682), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3270), .O(n3267), .CO(n3268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i23  (.I0(n7684), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3272), .O(n3269), .CO(n3270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i22  (.I0(n7686), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3274), .O(n3271), .CO(n3272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i21  (.I0(n7688), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3276), .O(n3273), .CO(n3274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i20  (.I0(n7690), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n3278), .O(n3275), .CO(n3276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2636/i19  (.I0(n7692), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2920), .O(n3277), .CO(n3278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2636/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2636/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i32  (.I0(n7701), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3289), .O(n3287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i31  (.I0(n7703), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3291), .O(n3288), .CO(n3289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i30  (.I0(n7705), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3293), .O(n3290), .CO(n3291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i29  (.I0(n7707), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3295), .O(n3292), .CO(n3293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i28  (.I0(n7709), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3297), .O(n3294), .CO(n3295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i27  (.I0(n7711), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3299), .O(n3296), .CO(n3297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i26  (.I0(n7713), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3301), .O(n3298), .CO(n3299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i25  (.I0(n7715), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3303), .O(n3300), .CO(n3301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i24  (.I0(n7717), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3305), .O(n3302), .CO(n3303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i23  (.I0(n7719), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3307), .O(n3304), .CO(n3305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i22  (.I0(n7721), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3309), .O(n3306), .CO(n3307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2552/i21  (.I0(n7723), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2843), .O(n3308), .CO(n3309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2552/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2552/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i32  (.I0(n7725), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3312), .O(n3310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i31  (.I0(n7727), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3314), .O(n3311), .CO(n3312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i30  (.I0(n7729), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3316), .O(n3313), .CO(n3314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i29  (.I0(n7731), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3318), .O(n3315), .CO(n3316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i28  (.I0(n7733), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3320), .O(n3317), .CO(n3318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i27  (.I0(n7735), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3328), .O(n3319), .CO(n3320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i26  (.I0(n7742), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3330), .O(n3327), .CO(n3328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i25  (.I0(n7744), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3332), .O(n3329), .CO(n3330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i24  (.I0(n7746), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3334), .O(n3331), .CO(n3332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2466/i23  (.I0(n7748), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2789), .O(n3333), .CO(n3334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2466/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2466/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i32  (.I0(n7750), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3337), .O(n3335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i31  (.I0(n7752), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3339), .O(n3336), .CO(n3337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i30  (.I0(n7754), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3341), .O(n3338), .CO(n3339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i29  (.I0(n7756), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3343), .O(n3340), .CO(n3341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i28  (.I0(n7758), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3345), .O(n3342), .CO(n3343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i27  (.I0(n7760), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3347), .O(n3344), .CO(n3345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i26  (.I0(n7762), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3349), .O(n3346), .CO(n3347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2378/i25  (.I0(n7764), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2747), .O(n3348), .CO(n3349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2378/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2378/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i3  (.I0(n2820), .I1(1'b0), .CI(n3353), 
            .O(n3350), .CO(n3351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i2  (.I0(n2822), .I1(n7221), .CI(1'b0), 
            .O(n3352), .CO(n3353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i32  (.I0(n7811), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3397), .O(n3395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i31  (.I0(n7813), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3399), .O(n3396), .CO(n3397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i30  (.I0(n7815), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3401), .O(n3398), .CO(n3399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i29  (.I0(n7817), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3403), .O(n3400), .CO(n3401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i28  (.I0(n7819), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3405), .O(n3402), .CO(n3403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2288/i27  (.I0(n7821), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2719), .O(n3404), .CO(n3405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2288/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2288/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i32  (.I0(n7823), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3408), .O(n3406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i31  (.I0(n7825), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3410), .O(n3407), .CO(n3408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i30  (.I0(n7827), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3412), .O(n3409), .CO(n3410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2196/i29  (.I0(n7829), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2689), .O(n3411), .CO(n3412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2196/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2196/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i32  (.I0(n7831), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3415), .O(n3413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_24/add_2102/i31  (.I0(n7833), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n2657), .O(n3414), .CO(n3415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \u_black_pixel_avg/div_24/add_2102/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_24/add_2102/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i1  (.I0(\u_rgb2dvi/enc_0/acc[0] ), .I1(n3492), 
            .CI(1'b0), .O(n3464), .CO(n3465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i2  (.I0(n2829), .I1(n7221), .CI(n12212), 
            .O(n3468), .CO(n3469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i1  (.I0(\u_rgb2dvi/enc_1/acc[0] ), .I1(n3492), 
            .CI(1'b0), .O(n3478), .CO(n3479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i1  (.I0(\u_rgb2dvi/enc_2/acc[0] ), .I1(n3492), 
            .CI(1'b0), .O(n3490), .CO(n3491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(1'b0), .I1(1'b1), .CI(n12213), 
            .O(n3492), .CO(n12214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i32  (.I0(n8230), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .CI(n3820), .O(n3818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i31  (.I0(n8232), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .CI(n3822), .O(n3819), .CO(n3820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i30  (.I0(n8234), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3824), .O(n3821), .CO(n3822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i29  (.I0(n8236), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3826), .O(n3823), .CO(n3824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i28  (.I0(n8238), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3828), .O(n3825), .CO(n3826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i27  (.I0(n8240), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3830), .O(n3827), .CO(n3828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i26  (.I0(n8242), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3832), .O(n3829), .CO(n3830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i25  (.I0(n8244), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3834), .O(n3831), .CO(n3832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i24  (.I0(n8246), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3836), .O(n3833), .CO(n3834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i23  (.I0(n8248), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3838), .O(n3835), .CO(n3836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i22  (.I0(n8250), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3840), .O(n3837), .CO(n3838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i21  (.I0(n8252), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3842), .O(n3839), .CO(n3840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i20  (.I0(n8254), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3844), .O(n3841), .CO(n3842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i19  (.I0(n8256), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n3846), .O(n3843), .CO(n3844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i18  (.I0(n8258), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n3848), .O(n3845), .CO(n3846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2718/i17  (.I0(n8260), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .CI(n2284), .O(n3847), .CO(n3848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2718/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2718/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i32  (.I0(n8262), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .CI(n3851), .O(n3849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i31  (.I0(n8264), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3853), .O(n3850), .CO(n3851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i30  (.I0(n8266), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3855), .O(n3852), .CO(n3853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i29  (.I0(n8268), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3857), .O(n3854), .CO(n3855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i28  (.I0(n8270), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3859), .O(n3856), .CO(n3857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i27  (.I0(n8272), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3861), .O(n3858), .CO(n3859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i26  (.I0(n8274), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3863), .O(n3860), .CO(n3861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i25  (.I0(n8276), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3865), .O(n3862), .CO(n3863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i24  (.I0(n8278), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3867), .O(n3864), .CO(n3865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i23  (.I0(n8280), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3869), .O(n3866), .CO(n3867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i22  (.I0(n8282), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3871), .O(n3868), .CO(n3869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i21  (.I0(n8284), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3873), .O(n3870), .CO(n3871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i20  (.I0(n8286), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n3875), .O(n3872), .CO(n3873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2636/i19  (.I0(n8288), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .CI(n2264), .O(n3874), .CO(n3875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2636/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2636/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i32  (.I0(n8290), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .CI(n3878), .O(n3876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i31  (.I0(n8292), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3880), .O(n3877), .CO(n3878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i30  (.I0(n8294), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3882), .O(n3879), .CO(n3880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i29  (.I0(n8296), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3884), .O(n3881), .CO(n3882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i28  (.I0(n8298), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3886), .O(n3883), .CO(n3884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i27  (.I0(n8300), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3888), .O(n3885), .CO(n3886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i26  (.I0(n8302), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3890), .O(n3887), .CO(n3888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i25  (.I0(n8304), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3892), .O(n3889), .CO(n3890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i24  (.I0(n8306), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3894), .O(n3891), .CO(n3892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i23  (.I0(n8308), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3896), .O(n3893), .CO(n3894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i22  (.I0(n8310), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n3898), .O(n3895), .CO(n3896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2552/i21  (.I0(n8312), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .CI(n2242), .O(n3897), .CO(n3898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2552/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2552/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i32  (.I0(n8314), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .CI(n3901), .O(n3899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i31  (.I0(n8316), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3903), .O(n3900), .CO(n3901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i30  (.I0(n8318), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3905), .O(n3902), .CO(n3903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i29  (.I0(n8320), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3907), .O(n3904), .CO(n3905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i28  (.I0(n8322), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3909), .O(n3906), .CO(n3907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i27  (.I0(n8324), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3911), .O(n3908), .CO(n3909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i26  (.I0(n8326), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3913), .O(n3910), .CO(n3911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i25  (.I0(n8328), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3915), .O(n3912), .CO(n3913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i24  (.I0(n8330), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n3917), .O(n3914), .CO(n3915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2466/i23  (.I0(n8332), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .CI(n2218), .O(n3916), .CO(n3917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2466/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2466/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i32  (.I0(n8334), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .CI(n3920), .O(n3918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i31  (.I0(n8336), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3922), .O(n3919), .CO(n3920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i30  (.I0(n8338), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3924), .O(n3921), .CO(n3922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i29  (.I0(n8340), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3926), .O(n3923), .CO(n3924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i28  (.I0(n8342), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3928), .O(n3925), .CO(n3926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i27  (.I0(n8344), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3930), .O(n3927), .CO(n3928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i26  (.I0(n8346), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n3932), .O(n3929), .CO(n3930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2378/i25  (.I0(n8348), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .CI(n2192), .O(n3931), .CO(n3932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2378/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2378/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i32  (.I0(n8350), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .CI(n3935), .O(n3933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i31  (.I0(n8352), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3937), .O(n3934), .CO(n3935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i30  (.I0(n8354), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3939), .O(n3936), .CO(n3937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i29  (.I0(n8356), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3941), .O(n3938), .CO(n3939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i28  (.I0(n8358), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n3943), .O(n3940), .CO(n3941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2288/i27  (.I0(n8360), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .CI(n2164), .O(n3942), .CO(n3943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2288/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2288/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i32  (.I0(n8362), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .CI(n3946), .O(n3944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i31  (.I0(n8364), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3948), .O(n3945), .CO(n3946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i30  (.I0(n8366), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n3950), .O(n3947), .CO(n3948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2196/i29  (.I0(n8368), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .CI(n2134), .O(n3949), .CO(n3950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2196/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2196/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i32  (.I0(n8370), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .CI(n3953), .O(n3951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/div_23/add_2102/i31  (.I0(n8372), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .CI(n2102), .O(n3952), .CO(n3953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \u_black_pixel_avg/div_23/add_2102/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/div_23/add_2102/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \u_black_pixel_avg/add_8/i32  (.I0(\u_black_pixel_avg/y_sum[31] ), 
            .I1(1'b0), .CI(n3956), .O(n3954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i31  (.I0(\u_black_pixel_avg/y_sum[30] ), 
            .I1(1'b0), .CI(n3958), .O(n3955), .CO(n3956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i30  (.I0(\u_black_pixel_avg/y_sum[29] ), 
            .I1(1'b0), .CI(n3960), .O(n3957), .CO(n3958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i29  (.I0(\u_black_pixel_avg/y_sum[28] ), 
            .I1(1'b0), .CI(n3962), .O(n3959), .CO(n3960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i28  (.I0(\u_black_pixel_avg/y_sum[27] ), 
            .I1(1'b0), .CI(n3964), .O(n3961), .CO(n3962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i27  (.I0(\u_black_pixel_avg/y_sum[26] ), 
            .I1(1'b0), .CI(n3966), .O(n3963), .CO(n3964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i26  (.I0(\u_black_pixel_avg/y_sum[25] ), 
            .I1(1'b0), .CI(n3968), .O(n3965), .CO(n3966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i25  (.I0(\u_black_pixel_avg/y_sum[24] ), 
            .I1(1'b0), .CI(n3970), .O(n3967), .CO(n3968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i24  (.I0(\u_black_pixel_avg/y_sum[23] ), 
            .I1(1'b0), .CI(n3972), .O(n3969), .CO(n3970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i23  (.I0(\u_black_pixel_avg/y_sum[22] ), 
            .I1(1'b0), .CI(n3974), .O(n3971), .CO(n3972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i22  (.I0(\u_black_pixel_avg/y_sum[21] ), 
            .I1(1'b0), .CI(n3976), .O(n3973), .CO(n3974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i21  (.I0(\u_black_pixel_avg/y_sum[20] ), 
            .I1(1'b0), .CI(n3978), .O(n3975), .CO(n3976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i20  (.I0(\u_black_pixel_avg/y_sum[19] ), 
            .I1(1'b0), .CI(n3980), .O(n3977), .CO(n3978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i19  (.I0(\u_black_pixel_avg/y_sum[18] ), 
            .I1(1'b0), .CI(n3982), .O(n3979), .CO(n3980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i18  (.I0(\u_black_pixel_avg/y_sum[17] ), 
            .I1(1'b0), .CI(n3984), .O(n3981), .CO(n3982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i17  (.I0(\u_black_pixel_avg/y_sum[16] ), 
            .I1(1'b0), .CI(n3986), .O(n3983), .CO(n3984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i16  (.I0(\u_black_pixel_avg/y_sum[15] ), 
            .I1(1'b0), .CI(n3988), .O(n3985), .CO(n3986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i15  (.I0(\u_black_pixel_avg/y_sum[14] ), 
            .I1(1'b0), .CI(n3990), .O(n3987), .CO(n3988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i14  (.I0(\u_black_pixel_avg/y_sum[13] ), 
            .I1(1'b0), .CI(n3992), .O(n3989), .CO(n3990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i13  (.I0(\u_black_pixel_avg/y_sum[12] ), 
            .I1(1'b0), .CI(n3994), .O(n3991), .CO(n3992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i12  (.I0(\u_black_pixel_avg/y_sum[11] ), 
            .I1(\lcd_ypos[11] ), .CI(n3996), .O(n3993), .CO(n3994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i11  (.I0(\u_black_pixel_avg/y_sum[10] ), 
            .I1(\lcd_ypos[10] ), .CI(n3998), .O(n3995), .CO(n3996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i10  (.I0(\u_black_pixel_avg/y_sum[9] ), 
            .I1(\lcd_ypos[9] ), .CI(n4000), .O(n3997), .CO(n3998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i9  (.I0(\u_black_pixel_avg/y_sum[8] ), 
            .I1(\lcd_ypos[8] ), .CI(n4002), .O(n3999), .CO(n4000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i8  (.I0(\u_black_pixel_avg/y_sum[7] ), 
            .I1(\lcd_ypos[7] ), .CI(n4004), .O(n4001), .CO(n4002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i7  (.I0(\u_black_pixel_avg/y_sum[6] ), 
            .I1(\lcd_ypos[6] ), .CI(n4006), .O(n4003), .CO(n4004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i6  (.I0(\u_black_pixel_avg/y_sum[5] ), 
            .I1(\lcd_ypos[5] ), .CI(n4008), .O(n4005), .CO(n4006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i5  (.I0(\u_black_pixel_avg/y_sum[4] ), 
            .I1(\lcd_ypos[4] ), .CI(n4010), .O(n4007), .CO(n4008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i4  (.I0(\u_black_pixel_avg/y_sum[3] ), 
            .I1(\lcd_ypos[3] ), .CI(n4012), .O(n4009), .CO(n4010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i3  (.I0(\u_black_pixel_avg/y_sum[2] ), 
            .I1(\lcd_ypos[2] ), .CI(n4014), .O(n4011), .CO(n4012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_8/i2  (.I0(\u_black_pixel_avg/y_sum[1] ), 
            .I1(\lcd_ypos[1] ), .CI(n1717), .O(n4013), .CO(n4014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(38)
    defparam \u_black_pixel_avg/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_8/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i32  (.I0(\u_black_pixel_avg/x_sum[31] ), 
            .I1(1'b0), .CI(n4017), .O(n4015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i32 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i31  (.I0(\u_black_pixel_avg/x_sum[30] ), 
            .I1(1'b0), .CI(n4019), .O(n4016), .CO(n4017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i30  (.I0(\u_black_pixel_avg/x_sum[29] ), 
            .I1(1'b0), .CI(n4021), .O(n4018), .CO(n4019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i29  (.I0(\u_black_pixel_avg/x_sum[28] ), 
            .I1(1'b0), .CI(n4023), .O(n4020), .CO(n4021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i28  (.I0(\u_black_pixel_avg/x_sum[27] ), 
            .I1(1'b0), .CI(n4025), .O(n4022), .CO(n4023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i27  (.I0(\u_black_pixel_avg/x_sum[26] ), 
            .I1(1'b0), .CI(n4027), .O(n4024), .CO(n4025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i26  (.I0(\u_black_pixel_avg/x_sum[25] ), 
            .I1(1'b0), .CI(n4029), .O(n4026), .CO(n4027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i25  (.I0(\u_black_pixel_avg/x_sum[24] ), 
            .I1(1'b0), .CI(n4031), .O(n4028), .CO(n4029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i24  (.I0(\u_black_pixel_avg/x_sum[23] ), 
            .I1(1'b0), .CI(n4033), .O(n4030), .CO(n4031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i23  (.I0(\u_black_pixel_avg/x_sum[22] ), 
            .I1(1'b0), .CI(n4035), .O(n4032), .CO(n4033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i22  (.I0(\u_black_pixel_avg/x_sum[21] ), 
            .I1(1'b0), .CI(n4037), .O(n4034), .CO(n4035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i21  (.I0(\u_black_pixel_avg/x_sum[20] ), 
            .I1(1'b0), .CI(n4039), .O(n4036), .CO(n4037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i20  (.I0(\u_black_pixel_avg/x_sum[19] ), 
            .I1(1'b0), .CI(n4041), .O(n4038), .CO(n4039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i19  (.I0(\u_black_pixel_avg/x_sum[18] ), 
            .I1(1'b0), .CI(n4043), .O(n4040), .CO(n4041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i18  (.I0(\u_black_pixel_avg/x_sum[17] ), 
            .I1(1'b0), .CI(n4045), .O(n4042), .CO(n4043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i17  (.I0(\u_black_pixel_avg/x_sum[16] ), 
            .I1(1'b0), .CI(n4047), .O(n4044), .CO(n4045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i16  (.I0(\u_black_pixel_avg/x_sum[15] ), 
            .I1(1'b0), .CI(n4049), .O(n4046), .CO(n4047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i15  (.I0(\u_black_pixel_avg/x_sum[14] ), 
            .I1(1'b0), .CI(n4051), .O(n4048), .CO(n4049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i14  (.I0(\u_black_pixel_avg/x_sum[13] ), 
            .I1(1'b0), .CI(n4053), .O(n4050), .CO(n4051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i13  (.I0(\u_black_pixel_avg/x_sum[12] ), 
            .I1(1'b0), .CI(n4055), .O(n4052), .CO(n4053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i12  (.I0(\u_black_pixel_avg/x_sum[11] ), 
            .I1(\lcd_xpos[11] ), .CI(n4057), .O(n4054), .CO(n4055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i11  (.I0(\u_black_pixel_avg/x_sum[10] ), 
            .I1(\lcd_xpos[10] ), .CI(n4059), .O(n4056), .CO(n4057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i10  (.I0(\u_black_pixel_avg/x_sum[9] ), 
            .I1(\lcd_xpos[9] ), .CI(n4061), .O(n4058), .CO(n4059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i9  (.I0(\u_black_pixel_avg/x_sum[8] ), 
            .I1(\lcd_xpos[8] ), .CI(n4063), .O(n4060), .CO(n4061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i8  (.I0(\u_black_pixel_avg/x_sum[7] ), 
            .I1(\lcd_xpos[7] ), .CI(n4065), .O(n4062), .CO(n4063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i7  (.I0(\u_black_pixel_avg/x_sum[6] ), 
            .I1(\lcd_xpos[6] ), .CI(n4067), .O(n4064), .CO(n4065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i6  (.I0(\u_black_pixel_avg/x_sum[5] ), 
            .I1(\lcd_xpos[5] ), .CI(n4069), .O(n4066), .CO(n4067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i5  (.I0(\u_black_pixel_avg/x_sum[4] ), 
            .I1(\lcd_xpos[4] ), .CI(n4071), .O(n4068), .CO(n4069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i4  (.I0(\u_black_pixel_avg/x_sum[3] ), 
            .I1(\lcd_xpos[3] ), .CI(n4073), .O(n4070), .CO(n4071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i3  (.I0(\u_black_pixel_avg/x_sum[2] ), 
            .I1(\lcd_xpos[2] ), .CI(n4075), .O(n4072), .CO(n4073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_7/i2  (.I0(\u_black_pixel_avg/x_sum[1] ), 
            .I1(\lcd_xpos[1] ), .CI(n1715), .O(n4074), .CO(n4075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(37)
    defparam \u_black_pixel_avg/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i31  (.I0(\u_black_pixel_avg/black_pixel_count[31] ), 
            .I1(1'b0), .CI(n4078), .O(n4076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i31 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i30  (.I0(\u_black_pixel_avg/black_pixel_count[30] ), 
            .I1(1'b0), .CI(n4080), .O(n4077), .CO(n4078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i30 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i29  (.I0(\u_black_pixel_avg/black_pixel_count[29] ), 
            .I1(1'b0), .CI(n4082), .O(n4079), .CO(n4080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i29 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i28  (.I0(\u_black_pixel_avg/black_pixel_count[28] ), 
            .I1(1'b0), .CI(n4084), .O(n4081), .CO(n4082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i28 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i27  (.I0(\u_black_pixel_avg/black_pixel_count[27] ), 
            .I1(1'b0), .CI(n4086), .O(n4083), .CO(n4084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i27 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i26  (.I0(\u_black_pixel_avg/black_pixel_count[26] ), 
            .I1(1'b0), .CI(n4088), .O(n4085), .CO(n4086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i26 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i25  (.I0(\u_black_pixel_avg/black_pixel_count[25] ), 
            .I1(1'b0), .CI(n4090), .O(n4087), .CO(n4088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i25 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i24  (.I0(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I1(1'b0), .CI(n4092), .O(n4089), .CO(n4090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i24 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i23  (.I0(\u_black_pixel_avg/black_pixel_count[23] ), 
            .I1(1'b0), .CI(n4094), .O(n4091), .CO(n4092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i23 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i22  (.I0(\u_black_pixel_avg/black_pixel_count[22] ), 
            .I1(1'b0), .CI(n4096), .O(n4093), .CO(n4094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i22 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i21  (.I0(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I1(1'b0), .CI(n4098), .O(n4095), .CO(n4096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i21 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i20  (.I0(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I1(1'b0), .CI(n4100), .O(n4097), .CO(n4098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i20 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i19  (.I0(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I1(1'b0), .CI(n4102), .O(n4099), .CO(n4100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i19 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i18  (.I0(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I1(1'b0), .CI(n4104), .O(n4101), .CO(n4102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i18 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i17  (.I0(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I1(1'b0), .CI(n4106), .O(n4103), .CO(n4104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i17 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i16  (.I0(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I1(1'b0), .CI(n4108), .O(n4105), .CO(n4106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i16 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i15  (.I0(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I1(1'b0), .CI(n4110), .O(n4107), .CO(n4108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i15 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i14  (.I0(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I1(1'b0), .CI(n4112), .O(n4109), .CO(n4110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i14 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i13  (.I0(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I1(1'b0), .CI(n4114), .O(n4111), .CO(n4112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i13 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i12  (.I0(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I1(1'b0), .CI(n4116), .O(n4113), .CO(n4114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i12 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i11  (.I0(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I1(1'b0), .CI(n4118), .O(n4115), .CO(n4116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i11 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i10  (.I0(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I1(1'b0), .CI(n4120), .O(n4117), .CO(n4118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i10 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i9  (.I0(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I1(1'b0), .CI(n4122), .O(n4119), .CO(n4120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i9 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i8  (.I0(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I1(1'b0), .CI(n4124), .O(n4121), .CO(n4122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i8 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i7  (.I0(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I1(1'b0), .CI(n4126), .O(n4123), .CO(n4124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i7 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i6  (.I0(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I1(1'b0), .CI(n4128), .O(n4125), .CO(n4126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i6 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i5  (.I0(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I1(1'b0), .CI(n4130), .O(n4127), .CO(n4128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i5 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i4  (.I0(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I1(1'b0), .CI(n4132), .O(n4129), .CO(n4130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i4 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i3  (.I0(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I1(1'b0), .CI(n4134), .O(n4131), .CO(n4132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i3 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_black_pixel_avg/add_34/i2  (.I0(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I1(1'b0), .CI(n1680), .O(n4133), .CO(n4134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(39)
    defparam \u_black_pixel_avg/add_34/i2 .I0_POLARITY = 1'b1;
    defparam \u_black_pixel_avg/add_34/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i12  (.I0(\u_lcd_driver/vcnt[11] ), 
            .I1(1'b1), .CI(n4137), .O(n4135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i11  (.I0(\u_lcd_driver/vcnt[10] ), 
            .I1(1'b1), .CI(n4139), .O(n4136), .CO(n4137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i10  (.I0(\u_lcd_driver/vcnt[9] ), 
            .I1(1'b1), .CI(n4141), .O(n4138), .CO(n4139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i9  (.I0(\u_lcd_driver/vcnt[8] ), .I1(1'b1), 
            .CI(n4143), .O(n4140), .CO(n4141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i8  (.I0(\u_lcd_driver/vcnt[7] ), .I1(1'b1), 
            .CI(n4145), .O(n4142), .CO(n4143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i7  (.I0(\u_lcd_driver/vcnt[6] ), .I1(1'b1), 
            .CI(n4147), .O(n4144), .CO(n4145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i6  (.I0(\u_lcd_driver/vcnt[5] ), .I1(1'b1), 
            .CI(n4149), .O(n4146), .CO(n4147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i5  (.I0(\u_lcd_driver/vcnt[4] ), .I1(1'b0), 
            .CI(n4151), .O(n4148), .CO(n4149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i4  (.I0(\u_lcd_driver/vcnt[3] ), .I1(1'b0), 
            .CI(n4153), .O(n4150), .CO(n4151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i3  (.I0(\u_lcd_driver/vcnt[2] ), .I1(1'b1), 
            .CI(n4155), .O(n4152), .CO(n4153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_61/add_2/i2  (.I0(\u_lcd_driver/vcnt[1] ), .I1(1'b1), 
            .CI(n1663), .O(n4154), .CO(n4155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \u_lcd_driver/sub_61/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_61/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i12  (.I0(\u_lcd_driver/hcnt[11] ), 
            .I1(1'b1), .CI(n4158), .O(n4156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i11  (.I0(\u_lcd_driver/hcnt[10] ), 
            .I1(1'b1), .CI(n4160), .O(n4157), .CO(n4158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i10  (.I0(\u_lcd_driver/hcnt[9] ), 
            .I1(1'b1), .CI(n4162), .O(n4159), .CO(n4160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i9  (.I0(\u_lcd_driver/hcnt[8] ), .I1(1'b0), 
            .CI(n4164), .O(n4161), .CO(n4162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i8  (.I0(\u_lcd_driver/hcnt[7] ), .I1(1'b1), 
            .CI(n4166), .O(n4163), .CO(n4164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i7  (.I0(\u_lcd_driver/hcnt[6] ), .I1(1'b1), 
            .CI(n4168), .O(n4165), .CO(n4166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i6  (.I0(\u_lcd_driver/hcnt[5] ), .I1(1'b1), 
            .CI(n4170), .O(n4167), .CO(n4168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i5  (.I0(\u_lcd_driver/hcnt[4] ), .I1(1'b1), 
            .CI(n4172), .O(n4169), .CO(n4170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i4  (.I0(\u_lcd_driver/hcnt[3] ), .I1(1'b1), 
            .CI(n4174), .O(n4171), .CO(n4172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/sub_60/add_2/i3  (.I0(\u_lcd_driver/hcnt[2] ), .I1(1'b1), 
            .CI(n1658), .O(n4173), .CO(n4174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \u_lcd_driver/sub_60/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/sub_60/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i11  (.I0(\u_lcd_driver/vcnt[11] ), .I1(1'b0), 
            .CI(n4177), .O(n4175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i10  (.I0(\u_lcd_driver/vcnt[10] ), .I1(1'b0), 
            .CI(n4179), .O(n4176), .CO(n4177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i9  (.I0(\u_lcd_driver/vcnt[9] ), .I1(1'b0), 
            .CI(n4181), .O(n4178), .CO(n4179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i8  (.I0(\u_lcd_driver/vcnt[8] ), .I1(1'b0), 
            .CI(n4183), .O(n4180), .CO(n4181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i7  (.I0(\u_lcd_driver/vcnt[7] ), .I1(1'b0), 
            .CI(n4185), .O(n4182), .CO(n4183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i6  (.I0(\u_lcd_driver/vcnt[6] ), .I1(1'b0), 
            .CI(n4187), .O(n4184), .CO(n4185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i5  (.I0(\u_lcd_driver/vcnt[5] ), .I1(1'b0), 
            .CI(n4189), .O(n4186), .CO(n4187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i4  (.I0(\u_lcd_driver/vcnt[4] ), .I1(1'b0), 
            .CI(n4191), .O(n4188), .CO(n4189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i3  (.I0(\u_lcd_driver/vcnt[3] ), .I1(1'b0), 
            .CI(n4193), .O(n4190), .CO(n4191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_82/i2  (.I0(\u_lcd_driver/vcnt[2] ), .I1(1'b0), 
            .CI(n1654), .O(n4192), .CO(n4193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_82/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_82/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i11  (.I0(\u_lcd_driver/hcnt[11] ), .I1(1'b0), 
            .CI(n4196), .O(n4194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i10  (.I0(\u_lcd_driver/hcnt[10] ), .I1(1'b0), 
            .CI(n4198), .O(n4195), .CO(n4196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i9  (.I0(\u_lcd_driver/hcnt[9] ), .I1(1'b0), 
            .CI(n4200), .O(n4197), .CO(n4198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i8  (.I0(\u_lcd_driver/hcnt[8] ), .I1(1'b0), 
            .CI(n4202), .O(n4199), .CO(n4200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i7  (.I0(\u_lcd_driver/hcnt[7] ), .I1(1'b0), 
            .CI(n4204), .O(n4201), .CO(n4202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i6  (.I0(\u_lcd_driver/hcnt[6] ), .I1(1'b0), 
            .CI(n4206), .O(n4203), .CO(n4204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i5  (.I0(\u_lcd_driver/hcnt[5] ), .I1(1'b0), 
            .CI(n4208), .O(n4205), .CO(n4206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i4  (.I0(\u_lcd_driver/hcnt[4] ), .I1(1'b0), 
            .CI(n4210), .O(n4207), .CO(n4208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i3  (.I0(\u_lcd_driver/hcnt[3] ), .I1(1'b0), 
            .CI(n4212), .O(n4209), .CO(n4210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_77/i2  (.I0(\u_lcd_driver/hcnt[2] ), .I1(1'b0), 
            .CI(n1480), .O(n4211), .CO(n4212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_77/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_77/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i9  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .CI(n4222), .O(n4220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i8  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .CI(n4224), .O(n4221), .CO(n4222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i7  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .CI(n4226), .CO(n4224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i6  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .CI(n4228), .CO(n4226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i5  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .CI(n4230), .CO(n4228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i4  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .CI(n4232), .CO(n4230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i3  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] ), 
            .CI(n4234), .CO(n4232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i2  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] ), 
            .CI(n1225), .CO(n4234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1278)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_55/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i10  (.I0(1'b0), 
            .I1(1'b1), .CI(n4237), .O(n4235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i9  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .CI(n4239), .O(n4236), .CO(n4237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i8  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] ), .CI(n4241), 
            .O(n4238), .CO(n4239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i7  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] ), .CI(n4243), 
            .O(n4240), .CO(n4241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i6  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] ), .CI(n4245), 
            .O(n4242), .CO(n4243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i5  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] ), .CI(n4247), 
            .O(n4244), .CO(n4245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i4  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] ), .CI(n4249), 
            .O(n4246), .CO(n4247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i3  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] ), .CI(n4251), 
            .O(n4248), .CO(n4249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i2  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] ), .CI(n1209), 
            .O(n4250), .CO(n4251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i8  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I1(1'b0), .CI(n4254), .O(n4252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i7  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n4256), .O(n4253), .CO(n4254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i6  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n4258), .O(n4255), .CO(n4256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i5  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n4260), .O(n4257), .CO(n4258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i4  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n4262), .O(n4259), .CO(n4260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i3  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n4264), .O(n4261), .CO(n4262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i2  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n1206), .O(n4263), .CO(n4264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i8  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(1'b0), .CI(n4267), .O(n4265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i7  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n4269), .O(n4266), .CO(n4267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i6  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n4271), .O(n4268), .CO(n4269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i5  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n4273), .O(n4270), .CO(n4271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i4  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n4275), .O(n4272), .CO(n4273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i3  (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n1202), .O(n4274), .CO(n4275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/sub_131/add_2/i5  (.I0(\u_axi4_ctrl_0/rfifo_cnt[4] ), 
            .I1(1'b1), .CI(n4278), .O(n4276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(356)
    defparam \u_axi4_ctrl_0/sub_131/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/sub_131/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/sub_131/add_2/i4  (.I0(\u_axi4_ctrl_0/rfifo_cnt[3] ), 
            .I1(1'b1), .CI(n4280), .O(n4277), .CO(n4278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(356)
    defparam \u_axi4_ctrl_0/sub_131/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/sub_131/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/sub_131/add_2/i3  (.I0(\u_axi4_ctrl_0/rfifo_cnt[2] ), 
            .I1(1'b1), .CI(n4282), .O(n4279), .CO(n4280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(356)
    defparam \u_axi4_ctrl_0/sub_131/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/sub_131/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/sub_131/add_2/i2  (.I0(\u_axi4_ctrl_0/rfifo_cnt[1] ), 
            .I1(1'b1), .CI(n979), .O(n4281), .CO(n4282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(356)
    defparam \u_axi4_ctrl_0/sub_131/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/sub_131/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i9  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(n8651), .CI(n4285), .O(n4283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i8  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(n8654), .CI(n4287), .O(n4284), .CO(n4285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i7  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(n8657), .CI(n4289), .O(n4286), .CO(n4287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i6  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(n8660), .CI(n4291), .O(n4288), .CO(n4289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i5  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(n8663), .CI(n4292), .O(n4290), .CO(n4291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i4  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .I1(n8666), .CI(n4293), .CO(n4292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i3  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] ), 
            .I1(n8669), .CI(n4294), .CO(n4293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i2  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] ), 
            .I1(n8672), .CI(n977), .CO(n4294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i10  (.I0(1'b0), 
            .I1(1'b1), .CI(n4297), .O(n4295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i9  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .CI(n4299), .O(n4296), .CO(n4297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i8  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] ), .CI(n4301), 
            .O(n4298), .CO(n4299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i7  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] ), .CI(n4303), 
            .O(n4300), .CO(n4301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i6  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] ), .CI(n4305), 
            .O(n4302), .CO(n4303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i5  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] ), .CI(n4307), 
            .O(n4304), .CO(n4305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i4  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] ), .CI(n4309), 
            .O(n4306), .CO(n4307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i3  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] ), .CI(n4311), 
            .O(n4308), .CO(n4309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i2  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] ), .CI(n962), 
            .O(n4310), .CO(n4311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i8  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I1(1'b0), .CI(n4314), .O(n4312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i7  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n4316), .O(n4313), .CO(n4314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i6  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n4318), .O(n4315), .CO(n4316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i5  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n4320), .O(n4317), .CO(n4318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i4  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n4322), .O(n4319), .CO(n4320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i3  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n4324), .O(n4321), .CO(n4322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i2  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n959), .O(n4323), .CO(n4324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1298)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_98/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i8  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(1'b0), .CI(n4327), .O(n4325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i7  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n4329), .O(n4326), .CO(n4327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i6  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n4331), .O(n4328), .CO(n4329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i5  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n4333), .O(n4330), .CO(n4331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i4  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n4335), .O(n4332), .CO(n4333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i3  (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n955), .O(n4334), .CO(n4335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1288)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/add_96/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i13  (.I0(\DdrCtrl_ARADDR_0[21] ), .I1(1'b0), 
            .CI(n4351), .O(n4349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i12  (.I0(\DdrCtrl_ARADDR_0[20] ), .I1(1'b0), 
            .CI(n4353), .O(n4350), .CO(n4351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i11  (.I0(\DdrCtrl_ARADDR_0[19] ), .I1(1'b0), 
            .CI(n4355), .O(n4352), .CO(n4353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i10  (.I0(\DdrCtrl_ARADDR_0[18] ), .I1(1'b0), 
            .CI(n4357), .O(n4354), .CO(n4355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i9  (.I0(\DdrCtrl_ARADDR_0[17] ), .I1(1'b0), 
            .CI(n4359), .O(n4356), .CO(n4357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i8  (.I0(\DdrCtrl_ARADDR_0[16] ), .I1(1'b0), 
            .CI(n4361), .O(n4358), .CO(n4359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i7  (.I0(\DdrCtrl_ARADDR_0[15] ), .I1(1'b0), 
            .CI(n4363), .O(n4360), .CO(n4361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i6  (.I0(\DdrCtrl_ARADDR_0[14] ), .I1(1'b0), 
            .CI(n4365), .O(n4362), .CO(n4363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i5  (.I0(\DdrCtrl_ARADDR_0[13] ), .I1(1'b0), 
            .CI(n4367), .O(n4364), .CO(n4365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i4  (.I0(\DdrCtrl_ARADDR_0[12] ), .I1(1'b0), 
            .CI(n4369), .O(n4366), .CO(n4367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_420/i3  (.I0(\DdrCtrl_ARADDR_0[11] ), .I1(1'b0), 
            .CI(n632), .O(n4368), .CO(n4369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(563)
    defparam \u_axi4_ctrl_0/add_420/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_420/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i8  (.I0(\u_axi4_ctrl_0/rc_burst[7] ), .I1(1'b0), 
            .CI(n4372), .O(n4370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i7  (.I0(\u_axi4_ctrl_0/rc_burst[6] ), .I1(1'b0), 
            .CI(n4374), .O(n4371), .CO(n4372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i6  (.I0(\u_axi4_ctrl_0/rc_burst[5] ), .I1(1'b0), 
            .CI(n4376), .O(n4373), .CO(n4374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i5  (.I0(\u_axi4_ctrl_0/rc_burst[4] ), .I1(1'b0), 
            .CI(n4378), .O(n4375), .CO(n4376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i4  (.I0(\u_axi4_ctrl_0/rc_burst[3] ), .I1(1'b0), 
            .CI(n4380), .O(n4377), .CO(n4378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i3  (.I0(\u_axi4_ctrl_0/rc_burst[2] ), .I1(1'b0), 
            .CI(n4382), .O(n4379), .CO(n4380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl_0/add_63/i2  (.I0(\u_axi4_ctrl_0/rc_burst[1] ), .I1(1'b0), 
            .CI(n547), .O(n4381), .CO(n4382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(251)
    defparam \u_axi4_ctrl_0/add_63/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/add_63/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i11  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[11] ), 
            .I1(1'b0), .CI(n4385), .O(n4383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i11 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i10  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[10] ), 
            .I1(1'b0), .CI(n4387), .O(n4384), .CO(n4385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i10 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i9  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[9] ), 
            .I1(1'b0), .CI(n4389), .O(n4386), .CO(n4387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i9 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i8  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[8] ), 
            .I1(1'b0), .CI(n4391), .O(n4388), .CO(n4389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i8 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i7  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[7] ), 
            .I1(1'b0), .CI(n4393), .O(n4390), .CO(n4391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i7 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i6  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[6] ), 
            .I1(1'b0), .CI(n4395), .O(n4392), .CO(n4393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i6 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i5  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[5] ), 
            .I1(1'b0), .CI(n4397), .O(n4394), .CO(n4395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i5 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i4  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[4] ), 
            .I1(1'b0), .CI(n4399), .O(n4396), .CO(n4397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i4 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i3  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[3] ), 
            .I1(1'b0), .CI(n4401), .O(n4398), .CO(n4399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i3 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_Sensor_Image_XYCrop_0/add_48/i2  (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[2] ), 
            .I1(1'b0), .CI(n542), .O(n4400), .CO(n4401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(94)
    defparam \u_Sensor_Image_XYCrop_0/add_48/i2 .I0_POLARITY = 1'b1;
    defparam \u_Sensor_Image_XYCrop_0/add_48/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i11  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[11] ), 
            .I1(1'b0), .CI(n4404), .O(n4402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i11 .I0_POLARITY = 1'b1;
    defparam \add_214/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i10  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[10] ), 
            .I1(1'b0), .CI(n4406), .O(n4403), .CO(n4404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i10 .I0_POLARITY = 1'b1;
    defparam \add_214/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i9  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[9] ), .I1(1'b0), 
            .CI(n4408), .O(n4405), .CO(n4406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i9 .I0_POLARITY = 1'b1;
    defparam \add_214/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i8  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[8] ), .I1(1'b0), 
            .CI(n4410), .O(n4407), .CO(n4408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i8 .I0_POLARITY = 1'b1;
    defparam \add_214/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i7  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[7] ), .I1(1'b0), 
            .CI(n4412), .O(n4409), .CO(n4410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i7 .I0_POLARITY = 1'b1;
    defparam \add_214/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i6  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[6] ), .I1(1'b0), 
            .CI(n4414), .O(n4411), .CO(n4412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i6 .I0_POLARITY = 1'b1;
    defparam \add_214/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i5  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[5] ), .I1(1'b0), 
            .CI(n4416), .O(n4413), .CO(n4414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i5 .I0_POLARITY = 1'b1;
    defparam \add_214/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i4  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[4] ), .I1(1'b0), 
            .CI(n4418), .O(n4415), .CO(n4416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i4 .I0_POLARITY = 1'b1;
    defparam \add_214/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i3  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[3] ), .I1(1'b0), 
            .CI(n4420), .O(n4417), .CO(n4418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i3 .I0_POLARITY = 1'b1;
    defparam \add_214/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_214/i2  (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[2] ), .I1(1'b0), 
            .CI(n464), .O(n4419), .CO(n4420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\Sensor_Image_XYCrop.v(113)
    defparam \add_214/i2 .I0_POLARITY = 1'b1;
    defparam \add_214/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i8  (.I0(\i2c_config_index[8] ), 
            .I1(1'b0), .CI(n4423), .O(n4421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i7  (.I0(\i2c_config_index[7] ), 
            .I1(1'b0), .CI(n4425), .O(n4422), .CO(n4423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i6  (.I0(\i2c_config_index[6] ), 
            .I1(1'b0), .CI(n4427), .O(n4424), .CO(n4425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i5  (.I0(\i2c_config_index[5] ), 
            .I1(1'b0), .CI(n4429), .O(n4426), .CO(n4427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i4  (.I0(\i2c_config_index[4] ), 
            .I1(1'b0), .CI(n4431), .O(n4428), .CO(n4429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i3  (.I0(\i2c_config_index[3] ), 
            .I1(1'b0), .CI(n4433), .O(n4430), .CO(n4431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_193/i2  (.I0(\i2c_config_index[2] ), 
            .I1(1'b0), .CI(n457), .O(n4432), .CO(n4433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(164)
    defparam \u_i2c_timing_ctrl_16bit/add_193/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_193/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i15  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[15] ), 
            .I1(1'b0), .CI(n4436), .O(n4434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i15 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i14  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[14] ), 
            .I1(1'b0), .CI(n4438), .O(n4435), .CO(n4436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i14 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i13  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[13] ), 
            .I1(1'b0), .CI(n4440), .O(n4437), .CO(n4438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i13 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i12  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[12] ), 
            .I1(1'b0), .CI(n4442), .O(n4439), .CO(n4440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i12 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i11  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[11] ), 
            .I1(1'b0), .CI(n4444), .O(n4441), .CO(n4442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i11 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i10  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[10] ), 
            .I1(1'b0), .CI(n4446), .O(n4443), .CO(n4444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i10 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i9  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[9] ), 
            .I1(1'b0), .CI(n4448), .O(n4445), .CO(n4446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i9 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i8  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[8] ), 
            .I1(1'b0), .CI(n4450), .O(n4447), .CO(n4448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i7  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[7] ), 
            .I1(1'b0), .CI(n4452), .O(n4449), .CO(n4450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i6  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[6] ), 
            .I1(1'b0), .CI(n4454), .O(n4451), .CO(n4452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i5  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[5] ), 
            .I1(1'b0), .CI(n4456), .O(n4453), .CO(n4454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i4  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[4] ), 
            .I1(1'b0), .CI(n4458), .O(n4455), .CO(n4456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i3  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[3] ), 
            .I1(1'b0), .CI(n4460), .O(n4457), .CO(n4458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_185/i2  (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[2] ), 
            .I1(1'b0), .CI(n454), .O(n4459), .CO(n4460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(102)
    defparam \u_i2c_timing_ctrl_16bit/add_185/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_185/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i26  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[26] ), 
            .I1(1'b0), .CI(n4463), .O(n4461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i26 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i25  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[25] ), 
            .I1(1'b0), .CI(n4465), .O(n4462), .CO(n4463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i25 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i24  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[24] ), 
            .I1(1'b0), .CI(n4467), .O(n4464), .CO(n4465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i24 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i23  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[23] ), 
            .I1(1'b0), .CI(n4469), .O(n4466), .CO(n4467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i23 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i22  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[22] ), 
            .I1(1'b0), .CI(n4471), .O(n4468), .CO(n4469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i22 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i21  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[21] ), 
            .I1(1'b0), .CI(n4473), .O(n4470), .CO(n4471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i21 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i20  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[20] ), 
            .I1(1'b0), .CI(n4475), .O(n4472), .CO(n4473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i20 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i19  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[19] ), 
            .I1(1'b0), .CI(n4477), .O(n4474), .CO(n4475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i19 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i18  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[18] ), 
            .I1(1'b0), .CI(n4479), .O(n4476), .CO(n4477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i18 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i17  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[17] ), 
            .I1(1'b0), .CI(n4481), .O(n4478), .CO(n4479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i17 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i16  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[16] ), 
            .I1(1'b0), .CI(n4483), .O(n4480), .CO(n4481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i16 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i15  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[15] ), 
            .I1(1'b0), .CI(n4485), .O(n4482), .CO(n4483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i15 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i14  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[14] ), 
            .I1(1'b0), .CI(n4487), .O(n4484), .CO(n4485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i14 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i13  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[13] ), 
            .I1(1'b0), .CI(n4489), .O(n4486), .CO(n4487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i13 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i12  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[12] ), 
            .I1(1'b0), .CI(n4491), .O(n4488), .CO(n4489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i12 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i11  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[11] ), 
            .I1(1'b0), .CI(n4493), .O(n4490), .CO(n4491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i11 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i10  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[10] ), 
            .I1(1'b0), .CI(n4495), .O(n4492), .CO(n4493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i10 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i9  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[9] ), 
            .I1(1'b0), .CI(n4497), .O(n4494), .CO(n4495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i9 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i8  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[8] ), 
            .I1(1'b0), .CI(n4499), .O(n4496), .CO(n4497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i7  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[7] ), 
            .I1(1'b0), .CI(n4501), .O(n4498), .CO(n4499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i6  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[6] ), 
            .I1(1'b0), .CI(n4503), .O(n4500), .CO(n4501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i5  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[5] ), 
            .I1(1'b0), .CI(n4505), .O(n4502), .CO(n4503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i4  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[4] ), 
            .I1(1'b0), .CI(n4507), .O(n4504), .CO(n4505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i3  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[3] ), 
            .I1(1'b0), .CI(n4509), .O(n4506), .CO(n4507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16bit/add_180/i2  (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[2] ), 
            .I1(1'b0), .CI(n432), .O(n4508), .CO(n4509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\cmos_i2c\i2c_timing_ctrl_16bit.v(67)
    defparam \u_i2c_timing_ctrl_16bit/add_180/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16bit/add_180/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), 
            .I1(1'b1), .CI(n4512), .O(n4510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I1(1'b1), .CI(n4514), .O(n4511), .CO(n4512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), 
            .I1(1'b1), .CI(n4516), .O(n4513), .CO(n4514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(1'b1), .CI(n4518), .O(n4515), .CO(n4516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), 
            .I1(1'b1), .CI(n4520), .O(n4517), .CO(n4518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I1(1'b1), .CI(n4522), .O(n4519), .CO(n4520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), 
            .I1(1'b1), .CI(n4524), .O(n4521), .CO(n4522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(1'b1), .CI(n4526), .O(n4523), .CO(n4524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), 
            .I1(1'b1), .CI(n4528), .O(n4525), .CO(n4526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I1(1'b1), .CI(n4530), .O(n4527), .CO(n4528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), 
            .I1(1'b1), .CI(n4532), .O(n4529), .CO(n4530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(1'b1), .CI(n4534), .O(n4531), .CO(n4532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), 
            .I1(1'b1), .CI(n4536), .O(n4533), .CO(n4534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I1(1'b1), .CI(n4538), .O(n4535), .CO(n4536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), 
            .I1(1'b1), .CI(n4540), .O(n4537), .CO(n4538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(1'b1), .CI(n4542), .O(n4539), .CO(n4540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), 
            .I1(1'b1), .CI(n4544), .O(n4541), .CO(n4542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I1(1'b1), .CI(n4546), .O(n4543), .CO(n4544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), 
            .I1(1'b1), .CI(n421), .O(n4545), .CO(n4546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i16  (.I0(n4566), .I1(n682), .CI(n4549), .O(n4547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i16 .I0_POLARITY = 1'b1;
    defparam \add_84/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i15  (.I0(n4567), .I1(n683), .CI(n4551), .O(n4548), 
            .CO(n4549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i15 .I0_POLARITY = 1'b1;
    defparam \add_84/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i14  (.I0(n4569), .I1(n684), .CI(n4553), .O(n4550), 
            .CO(n4551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i14 .I0_POLARITY = 1'b1;
    defparam \add_84/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i13  (.I0(n4571), .I1(n685), .CI(n4555), .O(n4552), 
            .CO(n4553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i13 .I0_POLARITY = 1'b1;
    defparam \add_84/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i12  (.I0(n4573), .I1(n686), .CI(n4557), .O(n4554), 
            .CO(n4555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i12 .I0_POLARITY = 1'b1;
    defparam \add_84/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i11  (.I0(n4575), .I1(n687), .CI(n4559), .O(n4556), 
            .CO(n4557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i11 .I0_POLARITY = 1'b1;
    defparam \add_84/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i10  (.I0(n4577), .I1(n688), .CI(n4561), .O(n4558), 
            .CO(n4559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i10 .I0_POLARITY = 1'b1;
    defparam \add_84/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i9  (.I0(n4579), .I1(n689), .CI(n4562), .O(n4560), 
            .CO(n4561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i9 .I0_POLARITY = 1'b1;
    defparam \add_84/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i8  (.I0(n4581), .I1(n690), .CI(n4563), .CO(n4562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i8 .I0_POLARITY = 1'b1;
    defparam \add_84/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i7  (.I0(n501), .I1(n691), .CI(n4564), .CO(n4563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i7 .I0_POLARITY = 1'b1;
    defparam \add_84/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i6  (.I0(n1649), .I1(n692), .CI(n4565), .CO(n4564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i6 .I0_POLARITY = 1'b1;
    defparam \add_84/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_84/i5  (.I0(n1651), .I1(n693), .CI(n419), .CO(n4565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_84/i5 .I0_POLARITY = 1'b1;
    defparam \add_84/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i16  (.I0(n617), .I1(n642), .CI(n4568), .O(n4566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i16 .I0_POLARITY = 1'b1;
    defparam \add_82/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i15  (.I0(n618), .I1(n643), .CI(n4570), .O(n4567), 
            .CO(n4568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i15 .I0_POLARITY = 1'b1;
    defparam \add_82/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i14  (.I0(n619), .I1(n644), .CI(n4572), .O(n4569), 
            .CO(n4570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i14 .I0_POLARITY = 1'b1;
    defparam \add_82/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i13  (.I0(n620), .I1(n8971), .CI(n4574), .O(n4571), 
            .CO(n4572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i13 .I0_POLARITY = 1'b1;
    defparam \add_82/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i12  (.I0(n621), .I1(n8974), .CI(n4576), .O(n4573), 
            .CO(n4574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i12 .I0_POLARITY = 1'b1;
    defparam \add_82/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i11  (.I0(n622), .I1(n647), .CI(n4578), .O(n4575), 
            .CO(n4576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i11 .I0_POLARITY = 1'b1;
    defparam \add_82/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i10  (.I0(n623), .I1(n648), .CI(n4580), .O(n4577), 
            .CO(n4578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i10 .I0_POLARITY = 1'b1;
    defparam \add_82/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i9  (.I0(n624), .I1(n649), .CI(n4582), .O(n4579), 
            .CO(n4580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i9 .I0_POLARITY = 1'b1;
    defparam \add_82/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_82/i8  (.I0(n625), .I1(n650), .CI(n502), .O(n4581), 
            .CO(n4582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam \add_82/i8 .I0_POLARITY = 1'b1;
    defparam \add_82/i8 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi0Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/r_wfifo_wdata[75] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[74] , \u_axi4_ctrl_0/r_wfifo_wdata[73] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[72] , \u_axi4_ctrl_0/r_wfifo_wdata[71] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[70] , \u_axi4_ctrl_0/r_wfifo_wdata[69] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[68] , \u_axi4_ctrl_0/r_wfifo_wdata[67] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[66] , \u_axi4_ctrl_0/r_wfifo_wdata[65] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[64] , \u_axi4_ctrl_0/r_wfifo_wdata[63] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[62] , \u_axi4_ctrl_0/r_wfifo_wdata[61] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[60] , \u_axi4_ctrl_0/r_wfifo_wdata[59] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[58] , \u_axi4_ctrl_0/r_wfifo_wdata[57] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[56] }), .WADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[67:48]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi0Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/r_wfifo_wdata[23] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[22] , \u_axi4_ctrl_0/r_wfifo_wdata[21] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[20] , \u_axi4_ctrl_0/r_wfifo_wdata[19] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[18] , \u_axi4_ctrl_0/r_wfifo_wdata[17] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[16] , \u_axi4_ctrl_0/r_wfifo_wdata[15] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[14] , \u_axi4_ctrl_0/r_wfifo_wdata[13] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[12] , \u_axi4_ctrl_0/r_wfifo_wdata[11] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[10] , \u_axi4_ctrl_0/r_wfifo_wdata[9] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[8] }), .WADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[15:0]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi0Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\r_XYCrop0_frame_Gray[7] , 
            \r_XYCrop0_frame_Gray[6] , \r_XYCrop0_frame_Gray[5] , \r_XYCrop0_frame_Gray[4] , 
            \r_XYCrop0_frame_Gray[3] , \r_XYCrop0_frame_Gray[2] , \r_XYCrop0_frame_Gray[1] , 
            \r_XYCrop0_frame_Gray[0] , \u_axi4_ctrl_0/r_wfifo_wdata[127] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[126] , \u_axi4_ctrl_0/r_wfifo_wdata[125] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[124] , \u_axi4_ctrl_0/r_wfifo_wdata[123] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[122] , \u_axi4_ctrl_0/r_wfifo_wdata[121] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[120] , \u_axi4_ctrl_0/r_wfifo_wdata[119] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[118] , \u_axi4_ctrl_0/r_wfifo_wdata[117] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[116] }), .WADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[127:108]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi0Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/r_wfifo_wdata[39] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[38] , \u_axi4_ctrl_0/r_wfifo_wdata[37] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[36] , \u_axi4_ctrl_0/r_wfifo_wdata[35] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[34] , \u_axi4_ctrl_0/r_wfifo_wdata[33] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[32] , \u_axi4_ctrl_0/r_wfifo_wdata[31] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[30] , \u_axi4_ctrl_0/r_wfifo_wdata[29] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[28] , \u_axi4_ctrl_0/r_wfifo_wdata[27] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[26] , \u_axi4_ctrl_0/r_wfifo_wdata[25] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[24] }), .WADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[31:16]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi0Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/r_wfifo_wdata[95] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[94] , \u_axi4_ctrl_0/r_wfifo_wdata[93] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[92] , \u_axi4_ctrl_0/r_wfifo_wdata[91] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[90] , \u_axi4_ctrl_0/r_wfifo_wdata[89] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[88] , \u_axi4_ctrl_0/r_wfifo_wdata[87] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[86] , \u_axi4_ctrl_0/r_wfifo_wdata[85] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[84] , \u_axi4_ctrl_0/r_wfifo_wdata[83] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[82] , \u_axi4_ctrl_0/r_wfifo_wdata[81] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[80] , \u_axi4_ctrl_0/r_wfifo_wdata[79] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[78] , \u_axi4_ctrl_0/r_wfifo_wdata[77] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[76] }), .WADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[87:68]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi0Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/r_wfifo_wdata[115] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[114] , \u_axi4_ctrl_0/r_wfifo_wdata[113] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[112] , \u_axi4_ctrl_0/r_wfifo_wdata[111] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[110] , \u_axi4_ctrl_0/r_wfifo_wdata[109] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[108] , \u_axi4_ctrl_0/r_wfifo_wdata[107] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[106] , \u_axi4_ctrl_0/r_wfifo_wdata[105] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[104] , \u_axi4_ctrl_0/r_wfifo_wdata[103] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[102] , \u_axi4_ctrl_0/r_wfifo_wdata[101] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[100] , \u_axi4_ctrl_0/r_wfifo_wdata[99] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[98] , \u_axi4_ctrl_0/r_wfifo_wdata[97] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[96] }), .WADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[107:88]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi0Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/r_wfifo_wdata[55] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[54] , \u_axi4_ctrl_0/r_wfifo_wdata[53] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[52] , \u_axi4_ctrl_0/r_wfifo_wdata[51] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[50] , \u_axi4_ctrl_0/r_wfifo_wdata[49] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[48] , \u_axi4_ctrl_0/r_wfifo_wdata[47] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[46] , \u_axi4_ctrl_0/r_wfifo_wdata[45] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[44] , \u_axi4_ctrl_0/r_wfifo_wdata[43] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[42] , \u_axi4_ctrl_0/r_wfifo_wdata[41] , 
            \u_axi4_ctrl_0/r_wfifo_wdata[40] }), .WADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[47:32]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\Axi0Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/rfifo_wdata[67] , 
            \u_axi4_ctrl_0/rfifo_wdata[66] , \u_axi4_ctrl_0/rfifo_wdata[65] , 
            \u_axi4_ctrl_0/rfifo_wdata[64] , \u_axi4_ctrl_0/rfifo_wdata[63] , 
            \u_axi4_ctrl_0/rfifo_wdata[62] , \u_axi4_ctrl_0/rfifo_wdata[61] , 
            \u_axi4_ctrl_0/rfifo_wdata[60] , \u_axi4_ctrl_0/rfifo_wdata[59] , 
            \u_axi4_ctrl_0/rfifo_wdata[58] , \u_axi4_ctrl_0/rfifo_wdata[57] , 
            \u_axi4_ctrl_0/rfifo_wdata[56] , \u_axi4_ctrl_0/rfifo_wdata[55] , 
            \u_axi4_ctrl_0/rfifo_wdata[54] , \u_axi4_ctrl_0/rfifo_wdata[53] , 
            \u_axi4_ctrl_0/rfifo_wdata[52] , \u_axi4_ctrl_0/rfifo_wdata[51] , 
            \u_axi4_ctrl_0/rfifo_wdata[50] , \u_axi4_ctrl_0/rfifo_wdata[49] , 
            \u_axi4_ctrl_0/rfifo_wdata[48] }), .WADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({\u_axi4_ctrl_0/w_rframe_data_gen[67] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[66] , \u_axi4_ctrl_0/w_rframe_data_gen[65] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[64] , \u_axi4_ctrl_0/w_rframe_data_gen[63] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[62] , \u_axi4_ctrl_0/w_rframe_data_gen[61] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[60] , \u_axi4_ctrl_0/w_rframe_data_gen[59] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[58] , \u_axi4_ctrl_0/w_rframe_data_gen[57] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[56] , \u_axi4_ctrl_0/w_rframe_data_gen[55] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[54] , \u_axi4_ctrl_0/w_rframe_data_gen[53] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[52] , \u_axi4_ctrl_0/w_rframe_data_gen[51] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[50] , \u_axi4_ctrl_0/w_rframe_data_gen[49] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[48] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\Axi0Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/rfifo_wdata[15] , 
            \u_axi4_ctrl_0/rfifo_wdata[14] , \u_axi4_ctrl_0/rfifo_wdata[13] , 
            \u_axi4_ctrl_0/rfifo_wdata[12] , \u_axi4_ctrl_0/rfifo_wdata[11] , 
            \u_axi4_ctrl_0/rfifo_wdata[10] , \u_axi4_ctrl_0/rfifo_wdata[9] , 
            \u_axi4_ctrl_0/rfifo_wdata[8] , \u_axi4_ctrl_0/rfifo_wdata[7] , 
            \u_axi4_ctrl_0/rfifo_wdata[6] , \u_axi4_ctrl_0/rfifo_wdata[5] , 
            \u_axi4_ctrl_0/rfifo_wdata[4] , \u_axi4_ctrl_0/rfifo_wdata[3] , 
            \u_axi4_ctrl_0/rfifo_wdata[2] , \u_axi4_ctrl_0/rfifo_wdata[1] , 
            \u_axi4_ctrl_0/rfifo_wdata[0] }), .WADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({\u_axi4_ctrl_0/w_rframe_data_gen[15] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[14] , \u_axi4_ctrl_0/w_rframe_data_gen[13] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[12] , \u_axi4_ctrl_0/w_rframe_data_gen[11] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[10] , \u_axi4_ctrl_0/w_rframe_data_gen[9] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[8] , \u_axi4_ctrl_0/w_rframe_data_gen[7] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[6] , \u_axi4_ctrl_0/w_rframe_data_gen[5] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[4] , \u_axi4_ctrl_0/w_rframe_data_gen[3] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[2] , \u_axi4_ctrl_0/w_rframe_data_gen[1] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1  (.WCLK(\Axi0Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/rfifo_wdata[127] , 
            \u_axi4_ctrl_0/rfifo_wdata[126] , \u_axi4_ctrl_0/rfifo_wdata[125] , 
            \u_axi4_ctrl_0/rfifo_wdata[124] , \u_axi4_ctrl_0/rfifo_wdata[123] , 
            \u_axi4_ctrl_0/rfifo_wdata[122] , \u_axi4_ctrl_0/rfifo_wdata[121] , 
            \u_axi4_ctrl_0/rfifo_wdata[120] , \u_axi4_ctrl_0/rfifo_wdata[119] , 
            \u_axi4_ctrl_0/rfifo_wdata[118] , \u_axi4_ctrl_0/rfifo_wdata[117] , 
            \u_axi4_ctrl_0/rfifo_wdata[116] , \u_axi4_ctrl_0/rfifo_wdata[115] , 
            \u_axi4_ctrl_0/rfifo_wdata[114] , \u_axi4_ctrl_0/rfifo_wdata[113] , 
            \u_axi4_ctrl_0/rfifo_wdata[112] , \u_axi4_ctrl_0/rfifo_wdata[111] , 
            \u_axi4_ctrl_0/rfifo_wdata[110] , \u_axi4_ctrl_0/rfifo_wdata[109] , 
            \u_axi4_ctrl_0/rfifo_wdata[108] }), .WADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({\u_axi4_ctrl_0/w_rframe_data_gen[127] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[126] , \u_axi4_ctrl_0/w_rframe_data_gen[125] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[124] , \u_axi4_ctrl_0/w_rframe_data_gen[123] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[122] , \u_axi4_ctrl_0/w_rframe_data_gen[121] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[120] , \u_axi4_ctrl_0/w_rframe_data_gen[119] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[118] , \u_axi4_ctrl_0/w_rframe_data_gen[117] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[116] , \u_axi4_ctrl_0/w_rframe_data_gen[115] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[114] , \u_axi4_ctrl_0/w_rframe_data_gen[113] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[112] , \u_axi4_ctrl_0/w_rframe_data_gen[111] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[110] , \u_axi4_ctrl_0/w_rframe_data_gen[109] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[108] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$f1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\Axi0Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/rfifo_wdata[31] , 
            \u_axi4_ctrl_0/rfifo_wdata[30] , \u_axi4_ctrl_0/rfifo_wdata[29] , 
            \u_axi4_ctrl_0/rfifo_wdata[28] , \u_axi4_ctrl_0/rfifo_wdata[27] , 
            \u_axi4_ctrl_0/rfifo_wdata[26] , \u_axi4_ctrl_0/rfifo_wdata[25] , 
            \u_axi4_ctrl_0/rfifo_wdata[24] , \u_axi4_ctrl_0/rfifo_wdata[23] , 
            \u_axi4_ctrl_0/rfifo_wdata[22] , \u_axi4_ctrl_0/rfifo_wdata[21] , 
            \u_axi4_ctrl_0/rfifo_wdata[20] , \u_axi4_ctrl_0/rfifo_wdata[19] , 
            \u_axi4_ctrl_0/rfifo_wdata[18] , \u_axi4_ctrl_0/rfifo_wdata[17] , 
            \u_axi4_ctrl_0/rfifo_wdata[16] }), .WADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({\u_axi4_ctrl_0/w_rframe_data_gen[31] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[30] , \u_axi4_ctrl_0/w_rframe_data_gen[29] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[28] , \u_axi4_ctrl_0/w_rframe_data_gen[27] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[26] , \u_axi4_ctrl_0/w_rframe_data_gen[25] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[24] , \u_axi4_ctrl_0/w_rframe_data_gen[23] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[22] , \u_axi4_ctrl_0/w_rframe_data_gen[21] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[20] , \u_axi4_ctrl_0/w_rframe_data_gen[19] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[18] , \u_axi4_ctrl_0/w_rframe_data_gen[17] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\Axi0Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/rfifo_wdata[87] , 
            \u_axi4_ctrl_0/rfifo_wdata[86] , \u_axi4_ctrl_0/rfifo_wdata[85] , 
            \u_axi4_ctrl_0/rfifo_wdata[84] , \u_axi4_ctrl_0/rfifo_wdata[83] , 
            \u_axi4_ctrl_0/rfifo_wdata[82] , \u_axi4_ctrl_0/rfifo_wdata[81] , 
            \u_axi4_ctrl_0/rfifo_wdata[80] , \u_axi4_ctrl_0/rfifo_wdata[79] , 
            \u_axi4_ctrl_0/rfifo_wdata[78] , \u_axi4_ctrl_0/rfifo_wdata[77] , 
            \u_axi4_ctrl_0/rfifo_wdata[76] , \u_axi4_ctrl_0/rfifo_wdata[75] , 
            \u_axi4_ctrl_0/rfifo_wdata[74] , \u_axi4_ctrl_0/rfifo_wdata[73] , 
            \u_axi4_ctrl_0/rfifo_wdata[72] , \u_axi4_ctrl_0/rfifo_wdata[71] , 
            \u_axi4_ctrl_0/rfifo_wdata[70] , \u_axi4_ctrl_0/rfifo_wdata[69] , 
            \u_axi4_ctrl_0/rfifo_wdata[68] }), .WADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({\u_axi4_ctrl_0/w_rframe_data_gen[87] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[86] , \u_axi4_ctrl_0/w_rframe_data_gen[85] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[84] , \u_axi4_ctrl_0/w_rframe_data_gen[83] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[82] , \u_axi4_ctrl_0/w_rframe_data_gen[81] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[80] , \u_axi4_ctrl_0/w_rframe_data_gen[79] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[78] , \u_axi4_ctrl_0/w_rframe_data_gen[77] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[76] , \u_axi4_ctrl_0/w_rframe_data_gen[75] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[74] , \u_axi4_ctrl_0/w_rframe_data_gen[73] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[72] , \u_axi4_ctrl_0/w_rframe_data_gen[71] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[70] , \u_axi4_ctrl_0/w_rframe_data_gen[69] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[68] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\Axi0Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/rfifo_wdata[107] , 
            \u_axi4_ctrl_0/rfifo_wdata[106] , \u_axi4_ctrl_0/rfifo_wdata[105] , 
            \u_axi4_ctrl_0/rfifo_wdata[104] , \u_axi4_ctrl_0/rfifo_wdata[103] , 
            \u_axi4_ctrl_0/rfifo_wdata[102] , \u_axi4_ctrl_0/rfifo_wdata[101] , 
            \u_axi4_ctrl_0/rfifo_wdata[100] , \u_axi4_ctrl_0/rfifo_wdata[99] , 
            \u_axi4_ctrl_0/rfifo_wdata[98] , \u_axi4_ctrl_0/rfifo_wdata[97] , 
            \u_axi4_ctrl_0/rfifo_wdata[96] , \u_axi4_ctrl_0/rfifo_wdata[95] , 
            \u_axi4_ctrl_0/rfifo_wdata[94] , \u_axi4_ctrl_0/rfifo_wdata[93] , 
            \u_axi4_ctrl_0/rfifo_wdata[92] , \u_axi4_ctrl_0/rfifo_wdata[91] , 
            \u_axi4_ctrl_0/rfifo_wdata[90] , \u_axi4_ctrl_0/rfifo_wdata[89] , 
            \u_axi4_ctrl_0/rfifo_wdata[88] }), .WADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({\u_axi4_ctrl_0/w_rframe_data_gen[107] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[106] , \u_axi4_ctrl_0/w_rframe_data_gen[105] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[104] , \u_axi4_ctrl_0/w_rframe_data_gen[103] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[102] , \u_axi4_ctrl_0/w_rframe_data_gen[101] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[100] , \u_axi4_ctrl_0/w_rframe_data_gen[99] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[98] , \u_axi4_ctrl_0/w_rframe_data_gen[97] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[96] , \u_axi4_ctrl_0/w_rframe_data_gen[95] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[94] , \u_axi4_ctrl_0/w_rframe_data_gen[93] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[92] , \u_axi4_ctrl_0/w_rframe_data_gen[91] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[90] , \u_axi4_ctrl_0/w_rframe_data_gen[89] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[88] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=20, WRITE_WIDTH=20, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 20;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\Axi0Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl_0/rfifo_wdata[47] , 
            \u_axi4_ctrl_0/rfifo_wdata[46] , \u_axi4_ctrl_0/rfifo_wdata[45] , 
            \u_axi4_ctrl_0/rfifo_wdata[44] , \u_axi4_ctrl_0/rfifo_wdata[43] , 
            \u_axi4_ctrl_0/rfifo_wdata[42] , \u_axi4_ctrl_0/rfifo_wdata[41] , 
            \u_axi4_ctrl_0/rfifo_wdata[40] , \u_axi4_ctrl_0/rfifo_wdata[39] , 
            \u_axi4_ctrl_0/rfifo_wdata[38] , \u_axi4_ctrl_0/rfifo_wdata[37] , 
            \u_axi4_ctrl_0/rfifo_wdata[36] , \u_axi4_ctrl_0/rfifo_wdata[35] , 
            \u_axi4_ctrl_0/rfifo_wdata[34] , \u_axi4_ctrl_0/rfifo_wdata[33] , 
            \u_axi4_ctrl_0/rfifo_wdata[32] }), .WADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] }), .RDATA({\u_axi4_ctrl_0/w_rframe_data_gen[47] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[46] , \u_axi4_ctrl_0/w_rframe_data_gen[45] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[44] , \u_axi4_ctrl_0/w_rframe_data_gen[43] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[42] , \u_axi4_ctrl_0/w_rframe_data_gen[41] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[40] , \u_axi4_ctrl_0/w_rframe_data_gen[39] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[38] , \u_axi4_ctrl_0/w_rframe_data_gen[37] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[36] , \u_axi4_ctrl_0/w_rframe_data_gen[35] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[34] , \u_axi4_ctrl_0/w_rframe_data_gen[33] , 
            \u_axi4_ctrl_0/w_rframe_data_gen[32] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(721)
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_MULT mult_80 (.CLK(\hdmi_clk1x_i~O ), .CEA(1'b1), .RSTA(1'b0), 
            .CEB(1'b0), .RSTB(1'b0), .CEO(1'b0), .RSTO(1'b0), .A({13'b0000000000000, 
            \u_axi4_ctrl_0/n1500 , \u_axi4_ctrl_0/n1501 , \u_axi4_ctrl_0/n1502 , 
            \u_axi4_ctrl_0/n1503 , \u_axi4_ctrl_0/n1504 }), .B({18'b000000000001001101}), 
            .O({Open_0, Open_1, Open_2, Open_3, Open_4, Open_5, 
            Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, 
            Open_13, Open_14, Open_15, Open_16, Open_17, Open_18, 
            Open_19, Open_20, Open_21, Open_22, n617, n618, n619, 
            n620, n621, n622, n623, n624, n625, n626, n627, 
            n628, n629})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b0, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b0, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam mult_80.WIDTH = 18;
    defparam mult_80.A_REG = 1'b1;
    defparam mult_80.B_REG = 1'b0;
    defparam mult_80.O_REG = 1'b0;
    defparam mult_80.CLK_POLARITY = 1'b1;
    defparam mult_80.CEA_POLARITY = 1'b1;
    defparam mult_80.RSTA_POLARITY = 1'b1;
    defparam mult_80.RSTA_SYNC = 1'b1;
    defparam mult_80.RSTA_VALUE = 1'b0;
    defparam mult_80.CEB_POLARITY = 1'b1;
    defparam mult_80.RSTB_POLARITY = 1'b1;
    defparam mult_80.RSTB_SYNC = 1'b0;
    defparam mult_80.RSTB_VALUE = 1'b0;
    defparam mult_80.CEO_POLARITY = 1'b1;
    defparam mult_80.RSTO_POLARITY = 1'b1;
    defparam mult_80.RSTO_SYNC = 1'b0;
    defparam mult_80.RSTO_VALUE = 1'b0;
    defparam mult_80.SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT mult_83 (.CLK(\hdmi_clk1x_i~O ), .CEA(1'b1), .RSTA(1'b0), 
            .CEB(1'b0), .RSTB(1'b0), .CEO(1'b0), .RSTO(1'b0), .A({13'b0000000000000, 
            \u_axi4_ctrl_0/n1495 , \u_axi4_ctrl_0/n1496 , \u_axi4_ctrl_0/n1497 , 
            \u_axi4_ctrl_0/n1498 , \u_axi4_ctrl_0/n1499 }), .B({18'b000000000000011101}), 
            .O({Open_23, Open_24, Open_25, Open_26, Open_27, Open_28, 
            Open_29, Open_30, Open_31, Open_32, Open_33, Open_34, 
            Open_35, Open_36, Open_37, Open_38, Open_39, Open_40, 
            Open_41, Open_42, Open_43, Open_44, Open_45, n682, n683, 
            n684, n685, n686, n687, n688, n689, n690, n691, 
            n692, n693, n694})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b0, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b0, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam mult_83.WIDTH = 18;
    defparam mult_83.A_REG = 1'b1;
    defparam mult_83.B_REG = 1'b0;
    defparam mult_83.O_REG = 1'b0;
    defparam mult_83.CLK_POLARITY = 1'b1;
    defparam mult_83.CEA_POLARITY = 1'b1;
    defparam mult_83.RSTA_POLARITY = 1'b1;
    defparam mult_83.RSTA_SYNC = 1'b1;
    defparam mult_83.RSTA_VALUE = 1'b0;
    defparam mult_83.CEB_POLARITY = 1'b1;
    defparam mult_83.RSTB_POLARITY = 1'b1;
    defparam mult_83.RSTB_SYNC = 1'b0;
    defparam mult_83.RSTB_VALUE = 1'b0;
    defparam mult_83.CEO_POLARITY = 1'b1;
    defparam mult_83.RSTO_POLARITY = 1'b1;
    defparam mult_83.RSTO_SYNC = 1'b0;
    defparam mult_83.RSTO_VALUE = 1'b0;
    defparam mult_83.SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT mult_81 (.CLK(\hdmi_clk1x_i~O ), .CEA(1'b1), .RSTA(1'b0), 
            .CEB(1'b0), .RSTB(1'b0), .CEO(1'b0), .RSTO(1'b0), .A({12'b000000000000, 
            \u_axi4_ctrl_0/n1505 , \u_axi4_ctrl_0/n1506 , \u_axi4_ctrl_0/n1507 , 
            \u_axi4_ctrl_0/n1492 , \u_axi4_ctrl_0/n1493 , \u_axi4_ctrl_0/n1494 }), 
            .B({18'b000000000001001011}), .O({Open_46, Open_47, Open_48, 
            Open_49, Open_50, Open_51, Open_52, Open_53, Open_54, 
            Open_55, Open_56, Open_57, Open_58, Open_59, Open_60, 
            Open_61, Open_62, Open_63, Open_64, Open_65, Open_66, 
            Open_67, Open_68, n642, n643, n644, n8971, n8974, 
            n647, n648, n649, n650, n651, n652, n653, n654})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b0, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b0, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\T35_Sensor_DDR3_LCD_Test.v(541)
    defparam mult_81.WIDTH = 18;
    defparam mult_81.A_REG = 1'b1;
    defparam mult_81.B_REG = 1'b0;
    defparam mult_81.O_REG = 1'b0;
    defparam mult_81.CLK_POLARITY = 1'b1;
    defparam mult_81.CEA_POLARITY = 1'b1;
    defparam mult_81.RSTA_POLARITY = 1'b1;
    defparam mult_81.RSTA_SYNC = 1'b1;
    defparam mult_81.RSTA_VALUE = 1'b0;
    defparam mult_81.CEB_POLARITY = 1'b1;
    defparam mult_81.RSTB_POLARITY = 1'b1;
    defparam mult_81.RSTB_SYNC = 1'b0;
    defparam mult_81.RSTB_VALUE = 1'b0;
    defparam mult_81.CEO_POLARITY = 1'b1;
    defparam mult_81.RSTO_POLARITY = 1'b1;
    defparam mult_81.RSTO_SYNC = 1'b0;
    defparam mult_81.RSTO_VALUE = 1'b0;
    defparam mult_81.SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__13703 (.I0(\DdrCtrl_ARADDR_0[21] ), .I1(\DdrCtrl_AWADDR_0[21] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13703.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13704 (.I0(\DdrCtrl_ARADDR_0[20] ), .I1(\DdrCtrl_AWADDR_0[20] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13704.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13705 (.I0(\DdrCtrl_ARADDR_0[19] ), .I1(\DdrCtrl_AWADDR_0[19] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13705.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13706 (.I0(\DdrCtrl_ARADDR_0[18] ), .I1(\DdrCtrl_AWADDR_0[18] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13706.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13707 (.I0(\DdrCtrl_ARADDR_0[17] ), .I1(\DdrCtrl_AWADDR_0[17] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13707.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13708 (.I0(\DdrCtrl_ARADDR_0[16] ), .I1(\DdrCtrl_AWADDR_0[16] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13708.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13709 (.I0(\DdrCtrl_ARADDR_0[15] ), .I1(\DdrCtrl_AWADDR_0[15] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13709.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13710 (.I0(\DdrCtrl_ARADDR_0[14] ), .I1(\DdrCtrl_AWADDR_0[14] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13710.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13711 (.I0(\DdrCtrl_ARADDR_0[13] ), .I1(\DdrCtrl_AWADDR_0[13] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13711.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13712 (.I0(\DdrCtrl_ARADDR_0[12] ), .I1(\DdrCtrl_AWADDR_0[12] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13712.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13713 (.I0(\DdrCtrl_ARADDR_0[11] ), .I1(\DdrCtrl_AWADDR_0[11] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13713.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13714 (.I0(\DdrCtrl_ARADDR_0[10] ), .I1(\DdrCtrl_AWADDR_0[10] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13714.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13715 (.I0(\DdrCtrl_ARADDR_0[9] ), .I1(\DdrCtrl_AWADDR_0[9] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13715.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13716 (.I0(\DdrCtrl_ARADDR_0[8] ), .I1(\DdrCtrl_AWADDR_0[8] ), 
            .I2(DdrCtrl_ATYPE_0), .O(DdrCtrl_AADDR_0[8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13716.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13717 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[7] ), 
            .O(DdrCtrl_AADDR_0[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13717.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13718 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[6] ), 
            .O(DdrCtrl_AADDR_0[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13718.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13719 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[5] ), 
            .O(DdrCtrl_AADDR_0[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13719.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13720 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[4] ), 
            .O(DdrCtrl_AADDR_0[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13720.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13721 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[3] ), 
            .O(DdrCtrl_AADDR_0[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13721.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13722 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[2] ), 
            .O(DdrCtrl_AADDR_0[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13722.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13723 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[1] ), 
            .O(DdrCtrl_AADDR_0[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13723.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13724 (.I0(DdrCtrl_ATYPE_0), .I1(\DdrCtrl_AWADDR_0[0] ), 
            .O(DdrCtrl_AADDR_0[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13724.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13725 (.I0(\u_axi4_ctrl_0/rc_burst[0] ), .I1(\u_axi4_ctrl_0/rc_burst[1] ), 
            .I2(\u_axi4_ctrl_0/rc_burst[2] ), .I3(\u_axi4_ctrl_0/rc_burst[3] ), 
            .O(n8988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13725.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13726 (.I0(\u_axi4_ctrl_0/rc_burst[4] ), .I1(\u_axi4_ctrl_0/rc_burst[5] ), 
            .I2(\u_axi4_ctrl_0/rc_burst[6] ), .I3(\u_axi4_ctrl_0/rc_burst[7] ), 
            .O(n8989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13726.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13727 (.I0(n8988), .I1(n8989), .O(DdrCtrl_WLAST_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__13727.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__13728 (.I0(\u_i2c_timing_ctrl_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16bit/current_state[2] ), .I2(\u_i2c_timing_ctrl_16bit/current_state[3] ), 
            .O(n8990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1e1e */ ;
    defparam LUT__13728.LUTMASK = 16'h1e1e;
    EFX_LUT4 LUT__13729 (.I0(\u_i2c_timing_ctrl_16bit/i2c_ctrl_clk ), .I1(n8990), 
            .O(cmos_sclk)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__13729.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__13730 (.I0(n8990), .I1(\u_i2c_timing_ctrl_16bit/current_state[0] ), 
            .O(cmos_sdat_OE)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__13730.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__13731 (.I0(\PowerOnResetCnt[4] ), .I1(\PowerOnResetCnt[5] ), 
            .I2(\PowerOnResetCnt[6] ), .I3(\PowerOnResetCnt[7] ), .O(n8991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13731.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13732 (.I0(\PowerOnResetCnt[0] ), .I1(\PowerOnResetCnt[1] ), 
            .I2(\PowerOnResetCnt[2] ), .I3(\PowerOnResetCnt[3] ), .O(n8992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13732.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13733 (.I0(n8991), .I1(n8992), .O(\reduce_nand_9/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13733.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13734 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), .O(n8993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13734.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13735 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), .O(n8994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13735.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13736 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), .O(n8995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13736.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13737 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), .O(n8996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13737.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13738 (.I0(n8993), .I1(n8994), .I2(n8995), .I3(n8996), 
            .O(n8997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13738.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13739 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), .O(n8998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13739.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13740 (.I0(n8997), .I1(n8998), .O(n8999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13740.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13741 (.I0(n8999), .I1(DdrInitDone), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__13741.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__13742 (.I0(\r_hdmi_tx0_o[7] ), .I1(\w_hdmi_txd0[0] ), 
            .I2(rc_hdmi_tx), .O(n927_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13742.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13743 (.I0(\r_hdmi_tx1_o[7] ), .I1(\w_hdmi_txd1[0] ), 
            .I2(rc_hdmi_tx), .O(n938_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13743.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13744 (.I0(\r_hdmi_tx2_o[7] ), .I1(\w_hdmi_txd2[0] ), 
            .I2(rc_hdmi_tx), .O(n949_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13744.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13745 (.I0(n1737), .I1(\PowerOnResetCnt[0] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n33_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__13745.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__13746 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .I2(DdrCtrl_CFG_SEQ_START), 
            .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__13746.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__13747 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__13747.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__13748 (.I0(n8999), .I1(n420), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13748.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13749 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__13749.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__13750 (.I0(n8999), .I1(n4545), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13750.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13751 (.I0(n8999), .I1(n4543), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13751.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13752 (.I0(n8999), .I1(n4541), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13752.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13753 (.I0(n8999), .I1(n4539), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13753.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13754 (.I0(n8999), .I1(n4537), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13754.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13755 (.I0(n8999), .I1(n4535), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13755.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13756 (.I0(n8999), .I1(n4533), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13756.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13757 (.I0(n8999), .I1(n4531), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13757.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13758 (.I0(n8999), .I1(n4529), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13758.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13759 (.I0(n8999), .I1(n4527), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13759.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13760 (.I0(n8999), .I1(n4525), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13760.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13761 (.I0(n8999), .I1(n4523), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13761.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13762 (.I0(n8999), .I1(n4521), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13762.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13763 (.I0(n8999), .I1(n4519), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13763.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13764 (.I0(n8999), .I1(n4517), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13764.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13765 (.I0(n8999), .I1(n4515), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13765.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13766 (.I0(n8999), .I1(n4513), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13766.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13767 (.I0(n8999), .I1(n4511), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13767.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13768 (.I0(n8999), .I1(n4510), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13768.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13769 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[0] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[1] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[2] ), .O(n9000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13769.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13770 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[4] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[5] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[6] ), .I3(\u_i2c_timing_ctrl_16bit/clk_cnt[7] ), 
            .O(n9001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13770.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13771 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[8] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[9] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[10] ), .O(n9002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13771.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13772 (.I0(n9000), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[3] ), 
            .I2(n9001), .I3(n9002), .O(n9003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__13772.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__13773 (.I0(n9003), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[11] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[12] ), .O(n9004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13773.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13774 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[19] ), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[25] ), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[18] ), .I3(\u_i2c_timing_ctrl_16bit/delay_cnt[26] ), 
            .O(n9005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13774.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13775 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[6] ), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[7] ), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[17] ), .I3(\u_i2c_timing_ctrl_16bit/delay_cnt[8] ), 
            .O(n9006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13775.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13776 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[9] ), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[10] ), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[11] ), .I3(\u_i2c_timing_ctrl_16bit/delay_cnt[12] ), 
            .O(n9007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13776.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13777 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[13] ), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[14] ), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[15] ), .I3(\u_i2c_timing_ctrl_16bit/delay_cnt[16] ), 
            .O(n9008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13777.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13778 (.I0(n9005), .I1(n9006), .I2(n9007), .I3(n9008), 
            .O(n9009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13778.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13779 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[20] ), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[21] ), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[22] ), .I3(\u_i2c_timing_ctrl_16bit/delay_cnt[23] ), 
            .O(n9010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13779.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13780 (.I0(n9010), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[24] ), 
            .O(n9011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13780.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13781 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[2] ), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[3] ), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[4] ), .I3(\u_i2c_timing_ctrl_16bit/delay_cnt[5] ), 
            .O(n9012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13781.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13782 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[1] ), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[0] ), 
            .I2(n9012), .O(n9013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13782.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13783 (.I0(n9009), .I1(n9011), .I2(n9013), .O(n9014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13783.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13784 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[14] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[15] ), 
            .I2(n9014), .O(n9015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13784.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13785 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[13] ), .I1(n9004), 
            .I2(n9015), .O(n9016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__13785.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__13786 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[0] ), .I1(n9016), 
            .O(\u_i2c_timing_ctrl_16bit/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13786.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13787 (.I0(\i2c_config_index[6] ), .I1(\i2c_config_index[7] ), 
            .O(n9017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13787.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13788 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .O(n9018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13788.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13789 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[5] ), 
            .O(n9019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13789.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13790 (.I0(n9018), .I1(n9019), .I2(n9017), .I3(\i2c_config_index[8] ), 
            .O(n9020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__13790.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__13791 (.I0(n9014), .I1(n9020), .I2(\u_i2c_timing_ctrl_16bit/current_state[0] ), 
            .I3(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), .O(n9021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf70f */ ;
    defparam LUT__13791.LUTMASK = 16'hf70f;
    EFX_LUT4 LUT__13792 (.I0(n9021), .I1(\u_i2c_timing_ctrl_16bit/current_state[1] ), 
            .I2(\u_i2c_timing_ctrl_16bit/current_state[2] ), .I3(\u_i2c_timing_ctrl_16bit/current_state[3] ), 
            .O(n9022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13792.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13793 (.I0(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] ), .I2(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3] ), .O(n9023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13793.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13794 (.I0(n9023), .I1(\u_i2c_timing_ctrl_16bit/current_state[0] ), 
            .I2(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), .I3(n8990), 
            .O(n9024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00 */ ;
    defparam LUT__13794.LUTMASK = 16'h2c00;
    EFX_LUT4 LUT__13795 (.I0(n9022), .I1(n9024), .O(n9025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13795.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13796 (.I0(\u_i2c_timing_ctrl_16bit/current_state[0] ), 
            .I1(n9025), .I2(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .O(\u_i2c_timing_ctrl_16bit/n189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__13796.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__13797 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[1] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[0] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[2] ), .I3(\u_i2c_timing_ctrl_16bit/clk_cnt[3] ), 
            .O(n9026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__13797.LUTMASK = 16'he000;
    EFX_LUT4 LUT__13798 (.I0(n9026), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[4] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[5] ), .I3(\u_i2c_timing_ctrl_16bit/clk_cnt[6] ), 
            .O(n9027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__13798.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__13799 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[7] ), .I1(n9027), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[8] ), .O(n9028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13799.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13800 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[9] ), .I1(n9028), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[10] ), .I3(\u_i2c_timing_ctrl_16bit/clk_cnt[11] ), 
            .O(n9029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__13800.LUTMASK = 16'he000;
    EFX_LUT4 LUT__13801 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[3] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[4] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[5] ), .O(n9030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13801.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13802 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[0] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[1] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[2] ), .I3(n9030), .O(n9031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__13802.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__13803 (.I0(n9031), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[6] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[7] ), .I3(\u_i2c_timing_ctrl_16bit/clk_cnt[8] ), 
            .O(n9032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13803.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13804 (.I0(n9032), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[9] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[10] ), .I3(\u_i2c_timing_ctrl_16bit/clk_cnt[11] ), 
            .O(n9033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__13804.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__13805 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[13] ), .I1(n9015), 
            .O(n9034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13805.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13806 (.I0(n9033), .I1(n9029), .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[12] ), 
            .I3(n9034), .O(\u_i2c_timing_ctrl_16bit/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__13806.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__13807 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[3] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[10] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[11] ), .I3(n9034), .O(n9035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13807.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13808 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[2] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[8] ), 
            .I2(\u_i2c_timing_ctrl_16bit/clk_cnt[9] ), .I3(\u_i2c_timing_ctrl_16bit/clk_cnt[12] ), 
            .O(n9036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13808.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13809 (.I0(\u_i2c_timing_ctrl_16bit/clk_cnt[0] ), .I1(\u_i2c_timing_ctrl_16bit/clk_cnt[1] ), 
            .I2(n9001), .I3(n9036), .O(n9037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13809.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13810 (.I0(n9035), .I1(n9037), .O(\u_i2c_timing_ctrl_16bit/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13810.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13814 (.I0(\u_i2c_timing_ctrl_16bit/current_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16bit/current_state[3] ), .O(n9040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13814.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13815 (.I0(\u_i2c_timing_ctrl_16bit/current_state[0] ), 
            .I1(n9040), .I2(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .I3(\u_i2c_timing_ctrl_16bit/current_state[1] ), .O(n9041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13815.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13816 (.I0(n9020), .I1(\i2c_config_index[0] ), .I2(n9041), 
            .O(\u_i2c_timing_ctrl_16bit/n241 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c2c */ ;
    defparam LUT__13816.LUTMASK = 16'h2c2c;
    EFX_LUT4 LUT__13817 (.I0(\u_i2c_timing_ctrl_16bit/current_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), .I2(\u_i2c_timing_ctrl_16bit/current_state[1] ), 
            .I3(n9040), .O(n9042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__13817.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__13818 (.I0(\u_i2c_timing_ctrl_16bit/current_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), .O(n9043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13818.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13819 (.I0(\u_i2c_timing_ctrl_16bit/current_state[3] ), 
            .I1(n9042), .I2(\u_i2c_timing_ctrl_16bit/current_state[1] ), 
            .I3(n9043), .O(n9044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcdd0 */ ;
    defparam LUT__13819.LUTMASK = 16'hcdd0;
    EFX_LUT4 LUT__13820 (.I0(n9043), .I1(\u_i2c_timing_ctrl_16bit/current_state[1] ), 
            .O(n9045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13820.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13821 (.I0(\u_i2c_timing_ctrl_16bit/current_state[3] ), 
            .I1(n9045), .I2(\u_i2c_timing_ctrl_16bit/current_state[2] ), 
            .O(n9046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__13821.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__13822 (.I0(n9044), .I1(n9046), .O(n9047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13822.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13823 (.I0(\u_i2c_timing_ctrl_16bit/current_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16bit/current_state[2] ), .I2(n9045), 
            .I3(n9042), .O(n9048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__13823.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__13824 (.I0(n9047), .I1(n9048), .O(n9049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13824.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13825 (.I0(n9044), .I1(n9048), .I2(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .O(n9050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__13825.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__13826 (.I0(n9049), .I1(n9025), .I2(n9050), .O(n9051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13826.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13827 (.I0(n9050), .I1(n9051), .I2(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), 
            .O(\u_i2c_timing_ctrl_16bit/n374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__13827.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__13828 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .O(n9052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13828.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13829 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .O(n9053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13829.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13830 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .O(n9054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13830.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13831 (.I0(n9052), .I1(n9053), .I2(n9054), .I3(\i2c_config_index[5] ), 
            .O(n9055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13831.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13832 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[3] ), 
            .O(n9056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13832.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13833 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[2] ), .O(n9057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h730d */ ;
    defparam LUT__13833.LUTMASK = 16'h730d;
    EFX_LUT4 LUT__13834 (.I0(\i2c_config_index[0] ), .I1(n9057), .I2(n9053), 
            .I3(n9056), .O(n9058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__13834.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__13835 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[5] ), 
            .O(n9059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13835.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13836 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .O(n9060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13836.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13837 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .O(n9061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13837.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13838 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[5] ), .I3(n9061), .O(n9062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__13838.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__13839 (.I0(\i2c_config_index[6] ), .I1(\i2c_config_index[7] ), 
            .O(n9063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13839.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13840 (.I0(n9060), .I1(n9059), .I2(n9062), .I3(n9063), 
            .O(n9064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__13840.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__13841 (.I0(n9055), .I1(n9058), .I2(\i2c_config_index[4] ), 
            .I3(n9064), .O(n9065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__13841.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__13842 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .O(n9066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13842.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13843 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[0] ), 
            .O(n9067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13843.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13844 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .O(n9068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13844.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13845 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .O(n9069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13845.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13846 (.I0(n9068), .I1(n9067), .I2(n9069), .O(n9070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13846.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13847 (.I0(\i2c_config_index[1] ), .I1(n9066), .I2(n9070), 
            .I3(\i2c_config_index[5] ), .O(n9071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__13847.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__13848 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .O(n9072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13848.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13849 (.I0(\i2c_config_index[0] ), .I1(n9072), .I2(n9054), 
            .O(n9073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__13849.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__13850 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[4] ), 
            .I2(n9073), .O(n9074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__13850.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__13851 (.I0(n9074), .I1(n9071), .I2(n9017), .O(n9075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13851.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13852 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[4] ), 
            .O(n9076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13852.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13853 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[2] ), .O(n9077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf6eb */ ;
    defparam LUT__13853.LUTMASK = 16'hf6eb;
    EFX_LUT4 LUT__13854 (.I0(n9052), .I1(n9076), .I2(n9077), .I3(\i2c_config_index[3] ), 
            .O(n9078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13854.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13855 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .O(n9079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13855.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13856 (.I0(n9079), .I1(\i2c_config_index[2] ), .I2(n9078), 
            .I3(\i2c_config_index[6] ), .O(n9080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd5f0 */ ;
    defparam LUT__13856.LUTMASK = 16'hd5f0;
    EFX_LUT4 LUT__13857 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[4] ), 
            .O(n9081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13857.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13858 (.I0(n9079), .I1(n9053), .I2(\i2c_config_index[2] ), 
            .I3(\i2c_config_index[6] ), .O(n9082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__13858.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__13859 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .O(n9083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13859.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13860 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[3] ), 
            .O(n9084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13860.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13861 (.I0(n9083), .I1(n9084), .I2(\i2c_config_index[4] ), 
            .O(n9085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__13861.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__13862 (.I0(n9085), .I1(n9082), .I2(n9052), .I3(\i2c_config_index[6] ), 
            .O(n9086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcafc */ ;
    defparam LUT__13862.LUTMASK = 16'hcafc;
    EFX_LUT4 LUT__13863 (.I0(\i2c_config_index[2] ), .I1(n9083), .O(n9087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13863.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13864 (.I0(n9018), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[4] ), .O(n9088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h070c */ ;
    defparam LUT__13864.LUTMASK = 16'h070c;
    EFX_LUT4 LUT__13865 (.I0(n9088), .I1(n9087), .I2(\i2c_config_index[6] ), 
            .I3(n9086), .O(n9089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__13865.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__13866 (.I0(n9081), .I1(n9067), .I2(\i2c_config_index[5] ), 
            .I3(n9089), .O(n9090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__13866.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__13867 (.I0(\i2c_config_index[5] ), .I1(n9080), .I2(n9090), 
            .I3(\i2c_config_index[7] ), .O(n9091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__13867.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__13868 (.I0(n9044), .I1(n9046), .O(n9092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13868.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13869 (.I0(n9075), .I1(n9091), .I2(n9065), .I3(n9092), 
            .O(n9093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__13869.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__13870 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[2] ), 
            .O(n9094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13870.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13871 (.I0(n9094), .I1(n9059), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[1] ), .O(n9095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he00f */ ;
    defparam LUT__13871.LUTMASK = 16'he00f;
    EFX_LUT4 LUT__13872 (.I0(\i2c_config_index[4] ), .I1(n9095), .I2(\i2c_config_index[5] ), 
            .I3(n9054), .O(n9096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030e */ ;
    defparam LUT__13872.LUTMASK = 16'h030e;
    EFX_LUT4 LUT__13873 (.I0(n9087), .I1(n9018), .I2(n9096), .I3(\i2c_config_index[4] ), 
            .O(n9097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__13873.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__13874 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[5] ), 
            .O(n9098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13874.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13875 (.I0(n9081), .I1(n9053), .I2(\i2c_config_index[3] ), 
            .I3(n9019), .O(n9099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__13875.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__13876 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[5] ), 
            .O(n9100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13876.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13877 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[3] ), 
            .O(n9101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13877.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13878 (.I0(n9100), .I1(n9101), .I2(n9098), .I3(n9099), 
            .O(n9102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__13878.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__13879 (.I0(n9095), .I1(n9102), .I2(n9097), .I3(\i2c_config_index[0] ), 
            .O(n9103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__13879.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__13880 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[4] ), 
            .O(n9104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13880.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13881 (.I0(n9104), .I1(n9066), .I2(\i2c_config_index[6] ), 
            .O(n9105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__13881.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__13882 (.I0(n9098), .I1(n9087), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[6] ), .O(n9106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__13882.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__13883 (.I0(n9105), .I1(n9103), .I2(n9106), .I3(\i2c_config_index[7] ), 
            .O(n9107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__13883.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__13884 (.I0(n9084), .I1(n9060), .O(n9108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13884.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13885 (.I0(\i2c_config_index[4] ), .I1(n9108), .I2(\i2c_config_index[5] ), 
            .O(n9109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__13885.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__13886 (.I0(n9109), .I1(\i2c_config_index[0] ), .I2(n9063), 
            .O(n9110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__13886.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__13887 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n9111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcb23 */ ;
    defparam LUT__13887.LUTMASK = 16'hcb23;
    EFX_LUT4 LUT__13888 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[3] ), .O(n9112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb35 */ ;
    defparam LUT__13888.LUTMASK = 16'heb35;
    EFX_LUT4 LUT__13889 (.I0(n9112), .I1(n9111), .I2(\i2c_config_index[4] ), 
            .O(n9113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__13889.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__13890 (.I0(\i2c_config_index[4] ), .I1(n9053), .I2(\i2c_config_index[3] ), 
            .I3(\i2c_config_index[0] ), .O(n9114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h45be */ ;
    defparam LUT__13890.LUTMASK = 16'h45be;
    EFX_LUT4 LUT__13891 (.I0(n9114), .I1(n9113), .I2(\i2c_config_index[5] ), 
            .I3(n9017), .O(n9115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__13891.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__13892 (.I0(n9107), .I1(n9110), .I2(n9115), .O(n9116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13892.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13893 (.I0(n9019), .I1(n9109), .I2(\i2c_config_index[6] ), 
            .O(n9117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__13893.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__13894 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[4] ), 
            .O(n9118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13894.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13895 (.I0(n9061), .I1(n9098), .I2(\i2c_config_index[3] ), 
            .O(n9119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13895.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13896 (.I0(\i2c_config_index[4] ), .I1(n9018), .I2(\i2c_config_index[1] ), 
            .I3(\i2c_config_index[5] ), .O(n9120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcfea */ ;
    defparam LUT__13896.LUTMASK = 16'hcfea;
    EFX_LUT4 LUT__13897 (.I0(n9083), .I1(n9067), .I2(n9119), .I3(n9120), 
            .O(n9121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__13897.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__13898 (.I0(n9118), .I1(n9017), .I2(n9121), .O(n9122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13898.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13899 (.I0(n9118), .I1(\i2c_config_index[3] ), .O(n9123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13899.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13900 (.I0(\i2c_config_index[5] ), .I1(n9123), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[1] ), .O(n9124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h68d7 */ ;
    defparam LUT__13900.LUTMASK = 16'h68d7;
    EFX_LUT4 LUT__13901 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[4] ), 
            .O(n9125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13901.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13902 (.I0(n9124), .I1(n9067), .I2(n9125), .I3(\i2c_config_index[3] ), 
            .O(n9126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__13902.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__13903 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[5] ), 
            .O(n9127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13903.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13904 (.I0(n9127), .I1(\i2c_config_index[4] ), .O(n9128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13904.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13905 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[2] ), 
            .O(n9129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13905.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13906 (.I0(n9098), .I1(n9128), .I2(\i2c_config_index[1] ), 
            .I3(n9129), .O(n9130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__13906.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__13907 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[4] ), .I3(n9018), .O(n9131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400 */ ;
    defparam LUT__13907.LUTMASK = 16'h1400;
    EFX_LUT4 LUT__13908 (.I0(n9130), .I1(n9131), .I2(\i2c_config_index[7] ), 
            .O(n9132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13908.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13909 (.I0(n9126), .I1(n9132), .I2(n9117), .I3(n9122), 
            .O(n9133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__13909.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__13910 (.I0(n9133), .I1(n9046), .I2(n9044), .I3(n9116), 
            .O(n9134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__13910.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__13911 (.I0(n9025), .I1(n9048), .I2(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .O(n9135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13911.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13912 (.I0(n9093), .I1(n9134), .I2(\u_i2c_timing_ctrl_16bit/i2c_wdata[0] ), 
            .I3(n9135), .O(n9136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__13912.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__13913 (.I0(n9049), .I1(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .O(n9137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13913.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13914 (.I0(n9136), .I1(n9137), .O(\u_i2c_timing_ctrl_16bit/n383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13914.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13922 (.I0(n9044), .I1(n9046), .O(n9143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13922.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13925 (.I0(n9046), .I1(n9044), .O(n9145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13925.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13931 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[8] ), .I1(n9007), 
            .I2(n9008), .I3(\u_i2c_timing_ctrl_16bit/delay_cnt[17] ), .O(n9149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__13931.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__13932 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[18] ), .I1(n9149), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[19] ), .O(n9150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__13932.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__13933 (.I0(n9150), .I1(n9011), .O(n9151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13933.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13934 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[25] ), .I1(n9151), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[26] ), .O(n9152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13934.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13935 (.I0(n431), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[1] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13935.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13936 (.I0(n9152), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[0] ), 
            .O(\u_i2c_timing_ctrl_16bit/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13936.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13937 (.I0(\u_i2c_timing_ctrl_16bit/i2c_wdata[3] ), .I1(\u_i2c_timing_ctrl_16bit/i2c_wdata[1] ), 
            .I2(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] ), 
            .O(n9153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__13937.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__13938 (.I0(\u_i2c_timing_ctrl_16bit/i2c_wdata[2] ), .I1(\u_i2c_timing_ctrl_16bit/i2c_wdata[0] ), 
            .I2(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] ), .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), 
            .O(n9154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__13938.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__13939 (.I0(\u_i2c_timing_ctrl_16bit/i2c_wdata[4] ), .I1(\u_i2c_timing_ctrl_16bit/i2c_wdata[6] ), 
            .I2(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] ), 
            .O(n9155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__13939.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__13940 (.I0(\u_i2c_timing_ctrl_16bit/i2c_wdata[5] ), .I1(\u_i2c_timing_ctrl_16bit/i2c_wdata[7] ), 
            .I2(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), .I3(n9155), 
            .O(n9156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__13940.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__13941 (.I0(n9154), .I1(n9153), .I2(n9156), .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2] ), 
            .O(n9157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__13941.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__13942 (.I0(n9157), .I1(n9049), .I2(n9050), .I3(n9025), 
            .O(n9158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__13942.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__13943 (.I0(n9024), .I1(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .I2(cmos_sdat_OUT), .I3(n9158), .O(\u_i2c_timing_ctrl_16bit/n369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__13943.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__13944 (.I0(n9016), .I1(n453), .O(\u_i2c_timing_ctrl_16bit/n157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13944.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13945 (.I0(n9016), .I1(n4459), .O(\u_i2c_timing_ctrl_16bit/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13945.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13946 (.I0(n9016), .I1(n4457), .O(\u_i2c_timing_ctrl_16bit/n155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13946.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13947 (.I0(n9016), .I1(n4455), .O(\u_i2c_timing_ctrl_16bit/n154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13947.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13948 (.I0(n9016), .I1(n4453), .O(\u_i2c_timing_ctrl_16bit/n153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13948.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13949 (.I0(n9016), .I1(n4451), .O(\u_i2c_timing_ctrl_16bit/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13949.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13950 (.I0(n9016), .I1(n4449), .O(\u_i2c_timing_ctrl_16bit/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13950.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13951 (.I0(n9016), .I1(n4447), .O(\u_i2c_timing_ctrl_16bit/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13951.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13952 (.I0(n9016), .I1(n4445), .O(\u_i2c_timing_ctrl_16bit/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13952.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13953 (.I0(n9016), .I1(n4443), .O(\u_i2c_timing_ctrl_16bit/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13953.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13954 (.I0(n9016), .I1(n4441), .O(\u_i2c_timing_ctrl_16bit/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13954.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13955 (.I0(n9016), .I1(n4439), .O(\u_i2c_timing_ctrl_16bit/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13955.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13956 (.I0(n9016), .I1(n4437), .O(\u_i2c_timing_ctrl_16bit/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13956.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13957 (.I0(n9016), .I1(n4435), .O(\u_i2c_timing_ctrl_16bit/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13957.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13958 (.I0(n9016), .I1(n4434), .O(\u_i2c_timing_ctrl_16bit/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13958.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13959 (.I0(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), .I1(\u_i2c_timing_ctrl_16bit/current_state[1] ), 
            .I2(n9044), .O(\u_i2c_timing_ctrl_16bit/n188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__13959.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__13960 (.I0(\u_i2c_timing_ctrl_16bit/current_state[2] ), 
            .I1(n9046), .I2(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .O(\u_i2c_timing_ctrl_16bit/n187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__13960.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__13961 (.I0(\u_i2c_timing_ctrl_16bit/current_state[3] ), 
            .I1(n9048), .I2(\u_i2c_timing_ctrl_16bit/i2c_transfer_en ), 
            .O(\u_i2c_timing_ctrl_16bit/n186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__13961.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__13962 (.I0(n456), .I1(n9020), .I2(\i2c_config_index[1] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__13962.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__13963 (.I0(n4432), .I1(n9020), .I2(\i2c_config_index[2] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n239 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13963.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13964 (.I0(n4430), .I1(n9020), .I2(\i2c_config_index[3] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13964.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13965 (.I0(n4428), .I1(n9020), .I2(\i2c_config_index[4] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n237 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13965.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13966 (.I0(n4426), .I1(n9020), .I2(\i2c_config_index[5] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13966.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13967 (.I0(n4424), .I1(n9020), .I2(\i2c_config_index[6] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13967.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13968 (.I0(n4422), .I1(n9020), .I2(\i2c_config_index[7] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__13968.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__13969 (.I0(n9020), .I1(n4421), .I2(\i2c_config_index[8] ), 
            .I3(n9041), .O(\u_i2c_timing_ctrl_16bit/n233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__13969.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__13970 (.I0(n9049), .I1(n9050), .I2(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), 
            .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] ), .O(\u_i2c_timing_ctrl_16bit/n373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__13970.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__13971 (.I0(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[1] ), .O(n9159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13971.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13972 (.I0(n9050), .I1(n9159), .I2(n9051), .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2] ), 
            .O(\u_i2c_timing_ctrl_16bit/n372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h75c0 */ ;
    defparam LUT__13972.LUTMASK = 16'h75c0;
    EFX_LUT4 LUT__13973 (.I0(n9159), .I1(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[2] ), 
            .O(n9160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13973.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13974 (.I0(n9050), .I1(n9160), .I2(n9051), .I3(\u_i2c_timing_ctrl_16bit/i2c_stream_cnt[3] ), 
            .O(\u_i2c_timing_ctrl_16bit/n371 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h75c0 */ ;
    defparam LUT__13974.LUTMASK = 16'h75c0;
    EFX_LUT4 LUT__13975 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[2] ), .O(n9161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfd4b */ ;
    defparam LUT__13975.LUTMASK = 16'hfd4b;
    EFX_LUT4 LUT__13976 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .O(n9162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__13976.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__13977 (.I0(n9162), .I1(n9161), .I2(\i2c_config_index[0] ), 
            .O(n9163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__13977.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__13978 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .O(n9164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13978.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13979 (.I0(n9061), .I1(n9094), .I2(n9164), .O(n9165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13979.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13980 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[0] ), .O(n9166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8baf */ ;
    defparam LUT__13980.LUTMASK = 16'h8baf;
    EFX_LUT4 LUT__13981 (.I0(n9166), .I1(n9165), .I2(\i2c_config_index[3] ), 
            .O(n9167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__13981.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__13982 (.I0(n9167), .I1(n9163), .I2(\i2c_config_index[5] ), 
            .I3(n9063), .O(n9168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__13982.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__13983 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .O(n9169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d3d */ ;
    defparam LUT__13983.LUTMASK = 16'h3d3d;
    EFX_LUT4 LUT__13984 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[0] ), .O(n9170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcbaf */ ;
    defparam LUT__13984.LUTMASK = 16'hcbaf;
    EFX_LUT4 LUT__13985 (.I0(n9170), .I1(n9169), .I2(\i2c_config_index[1] ), 
            .O(n9171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__13985.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__13986 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[0] ), .O(n9172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h775c */ ;
    defparam LUT__13986.LUTMASK = 16'h775c;
    EFX_LUT4 LUT__13987 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .O(n9173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13987.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13988 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[4] ), .O(n9174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6b6b */ ;
    defparam LUT__13988.LUTMASK = 16'h6b6b;
    EFX_LUT4 LUT__13989 (.I0(n9173), .I1(n9084), .I2(n9174), .O(n9175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__13989.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__13990 (.I0(n9171), .I1(n9172), .I2(n9175), .I3(\i2c_config_index[5] ), 
            .O(n9176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__13990.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__13991 (.I0(n9176), .I1(n9017), .I2(n9168), .I3(n9092), 
            .O(n9177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__13991.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__13992 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[5] ), .I3(\i2c_config_index[4] ), .O(n9178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c1f */ ;
    defparam LUT__13992.LUTMASK = 16'h2c1f;
    EFX_LUT4 LUT__13993 (.I0(n9056), .I1(n9104), .I2(\i2c_config_index[2] ), 
            .O(n9179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__13993.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__13994 (.I0(n9098), .I1(n9128), .I2(\i2c_config_index[1] ), 
            .I3(n9179), .O(n9180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__13994.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__13995 (.I0(\i2c_config_index[3] ), .I1(n9178), .I2(n9180), 
            .I3(\i2c_config_index[0] ), .O(n9181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__13995.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__13996 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[5] ), 
            .O(n9182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13996.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13997 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[1] ), 
            .O(n9183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13997.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13998 (.I0(n9100), .I1(n9066), .I2(n9052), .O(n9184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13998.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13999 (.I0(n9098), .I1(n9183), .I2(n9184), .I3(\i2c_config_index[6] ), 
            .O(n9185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__13999.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__14000 (.I0(n9131), .I1(n9182), .I2(\i2c_config_index[2] ), 
            .I3(n9185), .O(n9186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__14000.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__14001 (.I0(\i2c_config_index[3] ), .I1(n9053), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[4] ), .O(n9187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h233f */ ;
    defparam LUT__14001.LUTMASK = 16'h233f;
    EFX_LUT4 LUT__14002 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .O(n9188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14002.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14003 (.I0(n9084), .I1(n9083), .O(n9189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14003.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14004 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[2] ), 
            .O(n9190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14004.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14005 (.I0(\i2c_config_index[4] ), .I1(n9188), .I2(n9189), 
            .I3(n9190), .O(n9191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14005.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14006 (.I0(\i2c_config_index[2] ), .I1(n9052), .O(n9192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14006.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14007 (.I0(n9079), .I1(n9060), .I2(n9192), .I3(n9059), 
            .O(n9193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__14007.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__14008 (.I0(n9187), .I1(\i2c_config_index[5] ), .I2(n9191), 
            .I3(n9193), .O(n9194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14008.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14009 (.I0(n9183), .I1(n9190), .I2(n9173), .O(n9195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14009.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14010 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[5] ), 
            .O(n9196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14010.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14011 (.I0(n9060), .I1(n9196), .I2(n9094), .I3(\i2c_config_index[0] ), 
            .O(n9197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__14011.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__14012 (.I0(n9196), .I1(n9068), .I2(n9195), .I3(n9197), 
            .O(n9198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__14012.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__14013 (.I0(n9198), .I1(\i2c_config_index[3] ), .I2(\i2c_config_index[6] ), 
            .I3(n9194), .O(n9199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__14013.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__14014 (.I0(n9186), .I1(n9181), .I2(n9199), .I3(\i2c_config_index[7] ), 
            .O(n9200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__14014.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__14015 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .O(n9201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14015.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14016 (.I0(n9066), .I1(n9098), .I2(n9201), .O(n9202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14016.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14017 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[4] ), .O(n9203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h56e3 */ ;
    defparam LUT__14017.LUTMASK = 16'h56e3;
    EFX_LUT4 LUT__14018 (.I0(n9173), .I1(\i2c_config_index[3] ), .O(n9204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14018.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14019 (.I0(n9204), .I1(n9118), .I2(\i2c_config_index[1] ), 
            .O(n9205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d3d */ ;
    defparam LUT__14019.LUTMASK = 16'h3d3d;
    EFX_LUT4 LUT__14020 (.I0(\i2c_config_index[0] ), .I1(n9203), .I2(n9205), 
            .O(n9206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__14020.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__14021 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[4] ), .O(n9207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3 */ ;
    defparam LUT__14021.LUTMASK = 16'he3e3;
    EFX_LUT4 LUT__14022 (.I0(n9083), .I1(n9069), .I2(\i2c_config_index[0] ), 
            .I3(n9207), .O(n9208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40f */ ;
    defparam LUT__14022.LUTMASK = 16'hf40f;
    EFX_LUT4 LUT__14023 (.I0(n9208), .I1(n9206), .I2(\i2c_config_index[5] ), 
            .O(n9209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14023.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14024 (.I0(n9202), .I1(\i2c_config_index[1] ), .I2(n9209), 
            .I3(\i2c_config_index[6] ), .O(n9210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__14024.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__14025 (.I0(n9018), .I1(n9118), .I2(\i2c_config_index[0] ), 
            .O(n9211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14025.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14026 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .O(n9212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14026.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14027 (.I0(n9212), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[5] ), 
            .O(n9213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14027.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14028 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[2] ), 
            .O(n9214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14028.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14029 (.I0(n9070), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[4] ), .O(n9215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ca3 */ ;
    defparam LUT__14029.LUTMASK = 16'h3ca3;
    EFX_LUT4 LUT__14030 (.I0(\i2c_config_index[4] ), .I1(n9214), .I2(\i2c_config_index[5] ), 
            .I3(n9215), .O(n9216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__14030.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__14031 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[5] ), 
            .O(n9217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14031.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14032 (.I0(n9211), .I1(n9113), .I2(n9101), .I3(n9217), 
            .O(n9218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14032.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14033 (.I0(n9213), .I1(n9211), .I2(n9216), .I3(n9218), 
            .O(n9219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__14033.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__14034 (.I0(n9124), .I1(n9219), .I2(\i2c_config_index[6] ), 
            .O(n9220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14034.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14035 (.I0(n9220), .I1(n9210), .I2(n9044), .I3(\i2c_config_index[7] ), 
            .O(n9221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__14035.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__14036 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(n9214), .O(n9222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14036.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14037 (.I0(\i2c_config_index[1] ), .I1(n9067), .I2(n9222), 
            .I3(\i2c_config_index[4] ), .O(n9223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__14037.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__14038 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[1] ), .O(n9224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1554 */ ;
    defparam LUT__14038.LUTMASK = 16'h1554;
    EFX_LUT4 LUT__14039 (.I0(n9079), .I1(n9223), .I2(n9224), .I3(\i2c_config_index[5] ), 
            .O(n9225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__14039.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__14040 (.I0(n9087), .I1(n9098), .I2(n9225), .I3(\i2c_config_index[7] ), 
            .O(n9226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077 */ ;
    defparam LUT__14040.LUTMASK = 16'hf077;
    EFX_LUT4 LUT__14041 (.I0(n9196), .I1(n9066), .O(n9227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14041.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14042 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[4] ), 
            .O(n9228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14042.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14043 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[1] ), .O(n9229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h475f */ ;
    defparam LUT__14043.LUTMASK = 16'h475f;
    EFX_LUT4 LUT__14044 (.I0(n9069), .I1(n9228), .I2(n9229), .I3(\i2c_config_index[5] ), 
            .O(n9230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__14044.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__14045 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[3] ), .O(n9231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3002 */ ;
    defparam LUT__14045.LUTMASK = 16'h3002;
    EFX_LUT4 LUT__14046 (.I0(n9066), .I1(n9061), .I2(n9231), .I3(\i2c_config_index[1] ), 
            .O(n9232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__14046.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__14047 (.I0(n9123), .I1(n9230), .I2(n9232), .O(n9233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14047.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14048 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .O(n9234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14048.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14049 (.I0(n9234), .I1(\i2c_config_index[2] ), .I2(\i2c_config_index[3] ), 
            .I3(n9019), .O(n9235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__14049.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__14050 (.I0(n9227), .I1(n9233), .I2(n9235), .I3(\i2c_config_index[7] ), 
            .O(n9236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__14050.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__14051 (.I0(n9236), .I1(n9226), .I2(n9046), .I3(\i2c_config_index[6] ), 
            .O(n9237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__14051.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__14052 (.I0(n9200), .I1(n9177), .I2(n9221), .I3(n9237), 
            .O(n9238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__14052.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__14053 (.I0(\u_i2c_timing_ctrl_16bit/i2c_wdata[1] ), .I1(n9238), 
            .I2(n9137), .I3(n9135), .O(\u_i2c_timing_ctrl_16bit/n382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__14053.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__14054 (.I0(\i2c_config_index[0] ), .I1(n9056), .I2(\i2c_config_index[4] ), 
            .O(n9239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__14054.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__14055 (.I0(n9098), .I1(n9059), .I2(\i2c_config_index[0] ), 
            .O(n9240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14055.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14056 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[5] ), .O(n9241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fe8 */ ;
    defparam LUT__14056.LUTMASK = 16'h0fe8;
    EFX_LUT4 LUT__14057 (.I0(n9241), .I1(n9019), .I2(n9240), .I3(\i2c_config_index[2] ), 
            .O(n9242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd5f0 */ ;
    defparam LUT__14057.LUTMASK = 16'hd5f0;
    EFX_LUT4 LUT__14058 (.I0(\i2c_config_index[0] ), .I1(n9128), .I2(n9242), 
            .I3(\i2c_config_index[1] ), .O(n9243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcef0 */ ;
    defparam LUT__14058.LUTMASK = 16'hcef0;
    EFX_LUT4 LUT__14059 (.I0(n9239), .I1(n9113), .I2(\i2c_config_index[2] ), 
            .I3(n9243), .O(n9244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__14059.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__14060 (.I0(n9212), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[5] ), 
            .I3(\i2c_config_index[0] ), .O(n9245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h375f */ ;
    defparam LUT__14060.LUTMASK = 16'h375f;
    EFX_LUT4 LUT__14061 (.I0(n9212), .I1(\i2c_config_index[2] ), .I2(n9245), 
            .I3(n9063), .O(n9246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e00 */ ;
    defparam LUT__14061.LUTMASK = 16'h3e00;
    EFX_LUT4 LUT__14062 (.I0(n9079), .I1(\i2c_config_index[5] ), .I2(\i2c_config_index[6] ), 
            .O(n9247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__14062.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__14063 (.I0(\i2c_config_index[7] ), .I1(\i2c_config_index[6] ), 
            .O(n9248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14063.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14064 (.I0(n9247), .I1(n9201), .I2(n9164), .I3(n9248), 
            .O(n9249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__14064.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__14065 (.I0(n9076), .I1(n9247), .I2(\i2c_config_index[3] ), 
            .I3(n9201), .O(n9250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he300 */ ;
    defparam LUT__14065.LUTMASK = 16'he300;
    EFX_LUT4 LUT__14066 (.I0(n9060), .I1(n9087), .I2(n9247), .I3(\i2c_config_index[4] ), 
            .O(n9251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14066.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14067 (.I0(n9250), .I1(n9251), .O(n9252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14067.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14068 (.I0(n9125), .I1(n9101), .I2(\i2c_config_index[1] ), 
            .I3(\i2c_config_index[0] ), .O(n9253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h32f3 */ ;
    defparam LUT__14068.LUTMASK = 16'h32f3;
    EFX_LUT4 LUT__14069 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .O(n9254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14069.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14070 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .O(n9255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14070.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14071 (.I0(n9254), .I1(n9255), .I2(\i2c_config_index[5] ), 
            .O(n9256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14071.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14072 (.I0(\i2c_config_index[4] ), .I1(n9084), .I2(n9256), 
            .O(n9257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__14072.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__14073 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .O(n9258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14073.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14074 (.I0(n9258), .I1(n9127), .I2(\i2c_config_index[2] ), 
            .I3(n9052), .O(n9259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__14074.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__14075 (.I0(n9253), .I1(\i2c_config_index[2] ), .I2(n9257), 
            .I3(n9259), .O(n9260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__14075.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__14076 (.I0(\i2c_config_index[6] ), .I1(\i2c_config_index[7] ), 
            .O(n9261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14076.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14077 (.I0(n9252), .I1(n9260), .I2(n9261), .I3(n9249), 
            .O(n9262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__14077.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__14078 (.I0(n9017), .I1(n9244), .I2(n9246), .I3(n9262), 
            .O(n9263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__14078.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__14079 (.I0(n9182), .I1(n9234), .I2(\i2c_config_index[2] ), 
            .I3(\i2c_config_index[3] ), .O(n9264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa30 */ ;
    defparam LUT__14079.LUTMASK = 16'hfa30;
    EFX_LUT4 LUT__14080 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[1] ), .O(n9265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8aa2 */ ;
    defparam LUT__14080.LUTMASK = 16'h8aa2;
    EFX_LUT4 LUT__14081 (.I0(n9188), .I1(n9264), .I2(n9265), .O(n9266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14081.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14082 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[5] ), 
            .I2(\i2c_config_index[2] ), .I3(n9201), .O(n9267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8ee */ ;
    defparam LUT__14082.LUTMASK = 16'he8ee;
    EFX_LUT4 LUT__14083 (.I0(n9267), .I1(n9266), .I2(\i2c_config_index[4] ), 
            .I3(n9261), .O(n9268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__14083.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__14084 (.I0(n9127), .I1(n9060), .I2(n9268), .O(n9269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14084.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14085 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[2] ), .O(n9270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec57 */ ;
    defparam LUT__14085.LUTMASK = 16'hec57;
    EFX_LUT4 LUT__14086 (.I0(n9270), .I1(n9054), .I2(\i2c_config_index[4] ), 
            .O(n9271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__14086.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__14087 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[4] ), 
            .I2(n9129), .I3(n9059), .O(n9272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14087.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14088 (.I0(n9271), .I1(\i2c_config_index[5] ), .I2(n9272), 
            .I3(n9017), .O(n9273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__14088.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__14089 (.I0(n9109), .I1(n9235), .I2(n9063), .I3(n9046), 
            .O(n9274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__14089.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__14090 (.I0(n9269), .I1(n9273), .I2(n9274), .O(n9275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14090.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14091 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[3] ), .O(n9276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe4d */ ;
    defparam LUT__14091.LUTMASK = 16'hfe4d;
    EFX_LUT4 LUT__14092 (.I0(n9276), .I1(\i2c_config_index[4] ), .I2(\i2c_config_index[6] ), 
            .I3(\i2c_config_index[5] ), .O(n9277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfc0 */ ;
    defparam LUT__14092.LUTMASK = 16'hbfc0;
    EFX_LUT4 LUT__14093 (.I0(n9068), .I1(n9079), .I2(n9188), .I3(\i2c_config_index[5] ), 
            .O(n9278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__14093.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__14094 (.I0(n9067), .I1(n9255), .O(n9279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14094.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14095 (.I0(n9214), .I1(n9083), .I2(n9068), .O(n9280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__14095.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__14096 (.I0(n9279), .I1(n9167), .I2(\i2c_config_index[4] ), 
            .I3(n9280), .O(n9281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfca3 */ ;
    defparam LUT__14096.LUTMASK = 16'hfca3;
    EFX_LUT4 LUT__14097 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[3] ), 
            .O(n9282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14097.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14098 (.I0(n9060), .I1(n9282), .I2(n9129), .O(n9283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14098.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14099 (.I0(n9283), .I1(n9067), .I2(n9072), .I3(\i2c_config_index[4] ), 
            .O(n9284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3 */ ;
    defparam LUT__14099.LUTMASK = 16'haac3;
    EFX_LUT4 LUT__14100 (.I0(n9284), .I1(n9281), .I2(\i2c_config_index[5] ), 
            .O(n9285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__14100.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__14101 (.I0(n9278), .I1(n9129), .I2(n9285), .I3(\i2c_config_index[6] ), 
            .O(n9286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__14101.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__14102 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[2] ), .O(n9287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5cfb */ ;
    defparam LUT__14102.LUTMASK = 16'h5cfb;
    EFX_LUT4 LUT__14103 (.I0(n9287), .I1(n9286), .I2(\i2c_config_index[5] ), 
            .I3(n9277), .O(n9288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h35f3 */ ;
    defparam LUT__14103.LUTMASK = 16'h35f3;
    EFX_LUT4 LUT__14104 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[5] ), .O(n9289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff9 */ ;
    defparam LUT__14104.LUTMASK = 16'heff9;
    EFX_LUT4 LUT__14105 (.I0(n9094), .I1(n9127), .O(n9290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14105.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14106 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[5] ), .O(n9291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14106.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14107 (.I0(n9228), .I1(n9291), .I2(n9083), .O(n9292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14107.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14108 (.I0(n9234), .I1(n9290), .I2(n9292), .I3(\i2c_config_index[6] ), 
            .O(n9293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__14108.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__14109 (.I0(n9258), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[2] ), .O(n9294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001 */ ;
    defparam LUT__14109.LUTMASK = 16'h1001;
    EFX_LUT4 LUT__14110 (.I0(n9052), .I1(n9123), .I2(n9294), .I3(\i2c_config_index[5] ), 
            .O(n9295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__14110.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__14111 (.I0(n9061), .I1(\i2c_config_index[2] ), .I2(\i2c_config_index[1] ), 
            .I3(\i2c_config_index[3] ), .O(n9296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__14111.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__14112 (.I0(n9101), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[0] ), 
            .O(n9297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__14112.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__14113 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[0] ), .O(n9298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hba2f */ ;
    defparam LUT__14113.LUTMASK = 16'hba2f;
    EFX_LUT4 LUT__14114 (.I0(\i2c_config_index[3] ), .I1(n9061), .I2(\i2c_config_index[5] ), 
            .O(n9299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14114.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14115 (.I0(n9298), .I1(n9297), .I2(\i2c_config_index[2] ), 
            .I3(n9299), .O(n9300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__14115.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__14116 (.I0(n9296), .I1(n9295), .I2(n9300), .I3(\i2c_config_index[6] ), 
            .O(n9301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14116.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14117 (.I0(n9289), .I1(n9101), .I2(n9293), .I3(n9301), 
            .O(n9302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__14117.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__14118 (.I0(n9302), .I1(n9288), .I2(\i2c_config_index[7] ), 
            .I3(n9092), .O(n9303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__14118.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__14119 (.I0(n9044), .I1(n9263), .I2(n9275), .I3(n9303), 
            .O(n9304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__14119.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__14120 (.I0(\u_i2c_timing_ctrl_16bit/i2c_wdata[2] ), .I1(n9304), 
            .I2(n9137), .I3(n9135), .O(\u_i2c_timing_ctrl_16bit/n381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__14120.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__14121 (.I0(n9079), .I1(n9076), .I2(\i2c_config_index[5] ), 
            .O(n9305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14121.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14122 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[5] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[2] ), .O(n9306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3fe */ ;
    defparam LUT__14122.LUTMASK = 16'ha3fe;
    EFX_LUT4 LUT__14123 (.I0(n9231), .I1(\i2c_config_index[3] ), .I2(n9306), 
            .O(n9307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__14123.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__14124 (.I0(\i2c_config_index[0] ), .I1(n9305), .I2(n9307), 
            .O(n9308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__14124.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__14125 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[5] ), .O(n9309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7023 */ ;
    defparam LUT__14125.LUTMASK = 16'h7023;
    EFX_LUT4 LUT__14126 (.I0(n9309), .I1(n9019), .I2(\i2c_config_index[2] ), 
            .O(n9310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14126.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14127 (.I0(n9308), .I1(n9310), .I2(n9123), .I3(\i2c_config_index[1] ), 
            .O(n9311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec75 */ ;
    defparam LUT__14127.LUTMASK = 16'hec75;
    EFX_LUT4 LUT__14128 (.I0(n9130), .I1(\i2c_config_index[3] ), .I2(n9053), 
            .O(n9312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3 */ ;
    defparam LUT__14128.LUTMASK = 16'he3e3;
    EFX_LUT4 LUT__14129 (.I0(n9312), .I1(n9311), .I2(\i2c_config_index[6] ), 
            .O(n9313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__14129.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__14130 (.I0(n9018), .I1(\i2c_config_index[0] ), .I2(n9183), 
            .I3(n9196), .O(n9314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__14130.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__14131 (.I0(n9101), .I1(n9084), .I2(\i2c_config_index[1] ), 
            .O(n9315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14131.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14132 (.I0(n9072), .I1(n9228), .I2(n9315), .I3(n9190), 
            .O(n9316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__14132.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__14133 (.I0(\i2c_config_index[5] ), .I1(n9222), .I2(n9316), 
            .O(n9317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14133.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14134 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[1] ), .O(n9318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd73f */ ;
    defparam LUT__14134.LUTMASK = 16'hd73f;
    EFX_LUT4 LUT__14135 (.I0(n9234), .I1(\i2c_config_index[2] ), .I2(n9318), 
            .I3(\i2c_config_index[3] ), .O(n9319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__14135.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__14136 (.I0(n9062), .I1(\i2c_config_index[3] ), .I2(n9319), 
            .I3(\i2c_config_index[5] ), .O(n9320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf03b */ ;
    defparam LUT__14136.LUTMASK = 16'hf03b;
    EFX_LUT4 LUT__14137 (.I0(n9314), .I1(n9317), .I2(n9320), .I3(\i2c_config_index[6] ), 
            .O(n9321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__14137.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__14138 (.I0(n9321), .I1(n9313), .I2(\i2c_config_index[7] ), 
            .I3(n9143), .O(n9322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__14138.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__14139 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[5] ), 
            .I2(\i2c_config_index[2] ), .I3(n9079), .O(n9323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14139.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14140 (.I0(n9054), .I1(n9254), .I2(\i2c_config_index[4] ), 
            .I3(\i2c_config_index[5] ), .O(n9324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__14140.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__14141 (.I0(\i2c_config_index[3] ), .I1(n9076), .O(n9325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14141.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14142 (.I0(n9018), .I1(n9098), .I2(n9325), .I3(\i2c_config_index[1] ), 
            .O(n9326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__14142.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__14143 (.I0(n9098), .I1(\i2c_config_index[2] ), .I2(\i2c_config_index[3] ), 
            .O(n9327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__14143.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__14144 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[5] ), .O(n9328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdef3 */ ;
    defparam LUT__14144.LUTMASK = 16'hdef3;
    EFX_LUT4 LUT__14145 (.I0(n9328), .I1(n9327), .I2(\i2c_config_index[1] ), 
            .O(n9329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14145.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14146 (.I0(n9326), .I1(n9324), .I2(n9329), .I3(\i2c_config_index[0] ), 
            .O(n9330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__14146.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__14147 (.I0(n9104), .I1(n9188), .I2(n9067), .O(n9331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__14147.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__14148 (.I0(n9170), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[4] ), 
            .I3(\i2c_config_index[3] ), .O(n9332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcb00 */ ;
    defparam LUT__14148.LUTMASK = 16'hcb00;
    EFX_LUT4 LUT__14149 (.I0(\i2c_config_index[1] ), .I1(n9094), .I2(n9331), 
            .I3(n9332), .O(n9333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__14149.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__14150 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[2] ), 
            .I2(n9081), .O(n9334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__14150.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__14151 (.I0(n9118), .I1(n9334), .I2(n9084), .I3(\i2c_config_index[5] ), 
            .O(n9335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__14151.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__14152 (.I0(\i2c_config_index[5] ), .I1(n9333), .I2(n9335), 
            .O(n9336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14152.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14153 (.I0(n9330), .I1(n9323), .I2(n9336), .I3(\i2c_config_index[6] ), 
            .O(n9337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__14153.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__14154 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(n9053), .O(n9338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00 */ ;
    defparam LUT__14154.LUTMASK = 16'h2c00;
    EFX_LUT4 LUT__14155 (.I0(n9079), .I1(\i2c_config_index[1] ), .I2(n9123), 
            .I3(n9182), .O(n9339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__14155.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__14156 (.I0(\i2c_config_index[0] ), .I1(n9255), .I2(\i2c_config_index[4] ), 
            .I3(n9100), .O(n9340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__14156.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__14157 (.I0(n9339), .I1(n9340), .I2(n9017), .O(n9341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14157.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14158 (.I0(n9127), .I1(n9081), .I2(n9217), .O(n9342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14158.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14159 (.I0(n9254), .I1(\i2c_config_index[0] ), .I2(n9342), 
            .I3(n9018), .O(n9343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001 */ ;
    defparam LUT__14159.LUTMASK = 16'h1001;
    EFX_LUT4 LUT__14160 (.I0(n9127), .I1(n9087), .I2(\i2c_config_index[4] ), 
            .I3(\i2c_config_index[0] ), .O(n9344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__14160.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__14161 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[5] ), .I3(n9094), .O(n9345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc200 */ ;
    defparam LUT__14161.LUTMASK = 16'hc200;
    EFX_LUT4 LUT__14162 (.I0(\i2c_config_index[3] ), .I1(n9019), .I2(n9345), 
            .I3(n9063), .O(n9346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14162.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14163 (.I0(n9343), .I1(n9344), .I2(n9346), .O(n9347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14163.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14164 (.I0(n9338), .I1(\i2c_config_index[0] ), .I2(n9341), 
            .I3(n9347), .O(n9348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__14164.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__14165 (.I0(n9337), .I1(\i2c_config_index[7] ), .I2(n9348), 
            .I3(n9092), .O(n9349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__14165.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__14166 (.I0(n9166), .I1(n9078), .I2(\i2c_config_index[3] ), 
            .I3(\i2c_config_index[0] ), .O(n9350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5cc */ ;
    defparam LUT__14166.LUTMASK = 16'hc5cc;
    EFX_LUT4 LUT__14167 (.I0(n9118), .I1(n9188), .I2(\i2c_config_index[5] ), 
            .O(n9351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__14167.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__14168 (.I0(n9201), .I1(\i2c_config_index[2] ), .I2(\i2c_config_index[3] ), 
            .I3(n9019), .O(n9352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d00 */ ;
    defparam LUT__14168.LUTMASK = 16'h3d00;
    EFX_LUT4 LUT__14169 (.I0(n9351), .I1(n9352), .I2(\i2c_config_index[7] ), 
            .I3(n9350), .O(n9353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14169.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14170 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[3] ), .O(n9354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f */ ;
    defparam LUT__14170.LUTMASK = 16'hfe7f;
    EFX_LUT4 LUT__14171 (.I0(n9354), .I1(n9019), .I2(\i2c_config_index[7] ), 
            .O(n9355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__14171.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__14172 (.I0(n9054), .I1(n9087), .I2(\i2c_config_index[4] ), 
            .I3(\i2c_config_index[5] ), .O(n9356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfacf */ ;
    defparam LUT__14172.LUTMASK = 16'hfacf;
    EFX_LUT4 LUT__14173 (.I0(n9356), .I1(n9355), .I2(\i2c_config_index[6] ), 
            .I3(n9145), .O(n9357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__14173.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__14174 (.I0(n9353), .I1(n9357), .O(n9358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14174.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14175 (.I0(n9025), .I1(n9322), .I2(n9349), .I3(n9358), 
            .O(n9359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14175.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14176 (.I0(n9137), .I1(n9359), .I2(n9135), .I3(\u_i2c_timing_ctrl_16bit/i2c_wdata[3] ), 
            .O(\u_i2c_timing_ctrl_16bit/n380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcdc0 */ ;
    defparam LUT__14176.LUTMASK = 16'hcdc0;
    EFX_LUT4 LUT__14177 (.I0(n9188), .I1(\i2c_config_index[2] ), .I2(\i2c_config_index[4] ), 
            .O(n9360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__14177.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__14178 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[2] ), .O(n9361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h533f */ ;
    defparam LUT__14178.LUTMASK = 16'h533f;
    EFX_LUT4 LUT__14179 (.I0(n9094), .I1(n9052), .I2(\i2c_config_index[3] ), 
            .O(n9362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__14179.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__14180 (.I0(n9361), .I1(n9360), .I2(n9362), .I3(\i2c_config_index[0] ), 
            .O(n9363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__14180.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__14181 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[4] ), .O(n9364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h41f7 */ ;
    defparam LUT__14181.LUTMASK = 16'h41f7;
    EFX_LUT4 LUT__14182 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[1] ), .O(n9365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h35a3 */ ;
    defparam LUT__14182.LUTMASK = 16'h35a3;
    EFX_LUT4 LUT__14183 (.I0(n9365), .I1(n9364), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[5] ), .O(n9366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__14183.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__14184 (.I0(n9366), .I1(n9063), .O(n9367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14184.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14185 (.I0(n9079), .I1(n9248), .O(n9368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14185.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14186 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[5] ), .I3(\i2c_config_index[2] ), .O(n9369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb15 */ ;
    defparam LUT__14186.LUTMASK = 16'heb15;
    EFX_LUT4 LUT__14187 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[4] ), .O(n9370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd73c */ ;
    defparam LUT__14187.LUTMASK = 16'hd73c;
    EFX_LUT4 LUT__14188 (.I0(\i2c_config_index[3] ), .I1(n9183), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[4] ), .O(n9371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff3 */ ;
    defparam LUT__14188.LUTMASK = 16'heff3;
    EFX_LUT4 LUT__14189 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[4] ), .O(n9372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3 */ ;
    defparam LUT__14189.LUTMASK = 16'hedf3;
    EFX_LUT4 LUT__14190 (.I0(n9372), .I1(n9056), .I2(n9371), .I3(\i2c_config_index[5] ), 
            .O(n9373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__14190.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__14191 (.I0(n9370), .I1(n9059), .I2(n9373), .I3(n9017), 
            .O(n9374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__14191.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__14192 (.I0(n9369), .I1(n9368), .I2(n9374), .I3(n9092), 
            .O(n9375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14192.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14193 (.I0(n9363), .I1(\i2c_config_index[5] ), .I2(n9367), 
            .I3(n9375), .O(n9376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__14193.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__14194 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[5] ), .O(n9377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcc4 */ ;
    defparam LUT__14194.LUTMASK = 16'hfcc4;
    EFX_LUT4 LUT__14195 (.I0(n9127), .I1(\i2c_config_index[2] ), .I2(\i2c_config_index[4] ), 
            .I3(\i2c_config_index[1] ), .O(n9378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1c00 */ ;
    defparam LUT__14195.LUTMASK = 16'h1c00;
    EFX_LUT4 LUT__14196 (.I0(n9100), .I1(n9196), .I2(\i2c_config_index[1] ), 
            .I3(\i2c_config_index[3] ), .O(n9379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h35f3 */ ;
    defparam LUT__14196.LUTMASK = 16'h35f3;
    EFX_LUT4 LUT__14197 (.I0(\i2c_config_index[2] ), .I1(n9377), .I2(n9378), 
            .I3(n9379), .O(n9380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__14197.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__14198 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[5] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[3] ), .O(n9381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h75ea */ ;
    defparam LUT__14198.LUTMASK = 16'h75ea;
    EFX_LUT4 LUT__14199 (.I0(n9019), .I1(\i2c_config_index[2] ), .I2(n9381), 
            .I3(\i2c_config_index[1] ), .O(n9382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__14199.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__14200 (.I0(n9382), .I1(n9380), .I2(\i2c_config_index[0] ), 
            .O(n9383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14200.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14201 (.I0(n9098), .I1(n9214), .I2(n9383), .I3(n9261), 
            .O(n9384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__14201.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__14202 (.I0(n9190), .I1(n9068), .I2(n9212), .O(n9385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14202.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14203 (.I0(\i2c_config_index[2] ), .I1(n9019), .I2(n9189), 
            .I3(n9385), .O(n9386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__14203.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__14204 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[1] ), .O(n9387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030e */ ;
    defparam LUT__14204.LUTMASK = 16'h030e;
    EFX_LUT4 LUT__14205 (.I0(n9387), .I1(n9017), .I2(n9019), .O(n9388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14205.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14206 (.I0(n9386), .I1(n9261), .I2(n9388), .I3(n9145), 
            .O(n9389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__14206.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__14207 (.I0(n9087), .I1(\i2c_config_index[4] ), .I2(\i2c_config_index[6] ), 
            .O(n9390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__14207.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__14208 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[2] ), .O(n9391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h57ce */ ;
    defparam LUT__14208.LUTMASK = 16'h57ce;
    EFX_LUT4 LUT__14209 (.I0(n9391), .I1(\i2c_config_index[0] ), .I2(\i2c_config_index[3] ), 
            .I3(\i2c_config_index[5] ), .O(n9392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe00 */ ;
    defparam LUT__14209.LUTMASK = 16'hbe00;
    EFX_LUT4 LUT__14210 (.I0(n9201), .I1(\i2c_config_index[3] ), .I2(\i2c_config_index[2] ), 
            .I3(n9098), .O(n9393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b00 */ ;
    defparam LUT__14210.LUTMASK = 16'h4b00;
    EFX_LUT4 LUT__14211 (.I0(\i2c_config_index[2] ), .I1(n9255), .I2(n9392), 
            .I3(n9393), .O(n9394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__14211.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__14212 (.I0(n9119), .I1(\i2c_config_index[2] ), .I2(n9083), 
            .I3(n9125), .O(n9395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcb00 */ ;
    defparam LUT__14212.LUTMASK = 16'hcb00;
    EFX_LUT4 LUT__14213 (.I0(n9395), .I1(n9394), .I2(\i2c_config_index[6] ), 
            .I3(n9227), .O(n9396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__14213.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__14214 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[1] ), .O(n9397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf4d */ ;
    defparam LUT__14214.LUTMASK = 16'hbf4d;
    EFX_LUT4 LUT__14215 (.I0(n9228), .I1(\i2c_config_index[3] ), .I2(n9234), 
            .O(n9398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14215.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14216 (.I0(n9164), .I1(n9101), .I2(n9398), .I3(\i2c_config_index[5] ), 
            .O(n9399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__14216.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__14217 (.I0(n9397), .I1(n9059), .I2(n9399), .I3(n9017), 
            .O(n9400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__14217.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__14218 (.I0(n9108), .I1(\i2c_config_index[5] ), .I2(\i2c_config_index[4] ), 
            .I3(n9063), .O(n9401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__14218.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__14219 (.I0(n9400), .I1(n9401), .I2(n9143), .O(n9402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14219.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14220 (.I0(\i2c_config_index[7] ), .I1(n9396), .I2(n9390), 
            .I3(n9402), .O(n9403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__14220.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__14221 (.I0(n9384), .I1(n9376), .I2(n9389), .I3(n9403), 
            .O(n9404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__14221.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__14222 (.I0(n9137), .I1(\u_i2c_timing_ctrl_16bit/i2c_wdata[4] ), 
            .I2(n9404), .I3(n9135), .O(\u_i2c_timing_ctrl_16bit/n379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__14222.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__14223 (.I0(n9098), .I1(n9108), .I2(n9017), .O(n9405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__14223.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__14224 (.I0(n9084), .I1(n9387), .I2(n9019), .I3(n9405), 
            .O(n9406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__14224.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__14225 (.I0(n9083), .I1(\i2c_config_index[2] ), .I2(n9019), 
            .I3(n9385), .O(n9407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__14225.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__14226 (.I0(n9098), .I1(n9087), .I2(\i2c_config_index[6] ), 
            .I3(n9407), .O(n9408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__14226.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__14227 (.I0(n9408), .I1(\i2c_config_index[7] ), .O(n9409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14227.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14228 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[3] ), .O(n9410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2ff3 */ ;
    defparam LUT__14228.LUTMASK = 16'h2ff3;
    EFX_LUT4 LUT__14229 (.I0(n9279), .I1(n9222), .I2(n9410), .I3(\i2c_config_index[4] ), 
            .O(n9411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__14229.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__14230 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[1] ), .O(n9412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8ffe */ ;
    defparam LUT__14230.LUTMASK = 16'h8ffe;
    EFX_LUT4 LUT__14231 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[3] ), .O(n9413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'habb4 */ ;
    defparam LUT__14231.LUTMASK = 16'habb4;
    EFX_LUT4 LUT__14232 (.I0(n9413), .I1(n9412), .I2(\i2c_config_index[4] ), 
            .O(n9414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__14232.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__14233 (.I0(n9414), .I1(n9411), .I2(\i2c_config_index[5] ), 
            .O(n9415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__14233.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__14234 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(n9196), .I3(\i2c_config_index[3] ), .O(n9416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf5cf */ ;
    defparam LUT__14234.LUTMASK = 16'hf5cf;
    EFX_LUT4 LUT__14235 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[3] ), .I3(n9196), .O(n9417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1b2 */ ;
    defparam LUT__14235.LUTMASK = 16'he1b2;
    EFX_LUT4 LUT__14236 (.I0(n9417), .I1(n9416), .I2(\i2c_config_index[2] ), 
            .O(n9418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14236.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14237 (.I0(\i2c_config_index[5] ), .I1(n9234), .I2(n9079), 
            .I3(n9418), .O(n9419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef15 */ ;
    defparam LUT__14237.LUTMASK = 16'hef15;
    EFX_LUT4 LUT__14238 (.I0(n9415), .I1(n9419), .I2(\i2c_config_index[6] ), 
            .I3(\i2c_config_index[7] ), .O(n9420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__14238.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__14239 (.I0(\i2c_config_index[4] ), .I1(n9018), .I2(\i2c_config_index[0] ), 
            .I3(\i2c_config_index[5] ), .O(n9421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__14239.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__14240 (.I0(n9101), .I1(n9067), .I2(n9019), .I3(n9214), 
            .O(n9422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__14240.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__14241 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[3] ), .O(n9423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb0a */ ;
    defparam LUT__14241.LUTMASK = 16'heb0a;
    EFX_LUT4 LUT__14242 (.I0(\i2c_config_index[5] ), .I1(n9423), .I2(n9061), 
            .I3(n9214), .O(n9424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__14242.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__14243 (.I0(n9421), .I1(n9422), .I2(n9424), .I3(\i2c_config_index[1] ), 
            .O(n9425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__14243.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__14244 (.I0(\i2c_config_index[3] ), .I1(n9125), .I2(n9067), 
            .I3(n9425), .O(n9426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__14244.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__14245 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(n9079), .O(n9427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6100 */ ;
    defparam LUT__14245.LUTMASK = 16'h6100;
    EFX_LUT4 LUT__14246 (.I0(n9112), .I1(n9068), .I2(\i2c_config_index[3] ), 
            .I3(\i2c_config_index[4] ), .O(n9428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14246.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14247 (.I0(n9066), .I1(n9282), .I2(n9060), .O(n9429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__14247.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__14248 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[2] ), 
            .I2(n9188), .O(n9430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9e9e */ ;
    defparam LUT__14248.LUTMASK = 16'h9e9e;
    EFX_LUT4 LUT__14249 (.I0(n9430), .I1(n9429), .I2(\i2c_config_index[4] ), 
            .O(n9431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14249.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14250 (.I0(n9428), .I1(n9427), .I2(n9431), .I3(\i2c_config_index[5] ), 
            .O(n9432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__14250.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__14251 (.I0(n9426), .I1(n9432), .I2(\i2c_config_index[6] ), 
            .I3(n9420), .O(n9433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a */ ;
    defparam LUT__14251.LUTMASK = 16'hf30a;
    EFX_LUT4 LUT__14252 (.I0(n9409), .I1(n9406), .I2(n9433), .I3(n9046), 
            .O(n9434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__14252.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__14253 (.I0(n9228), .I1(n9162), .O(n9435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14253.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14254 (.I0(n9435), .I1(n9325), .I2(\i2c_config_index[5] ), 
            .I3(\i2c_config_index[0] ), .O(n9436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__14254.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__14255 (.I0(n9081), .I1(n9066), .I2(\i2c_config_index[5] ), 
            .I3(\i2c_config_index[7] ), .O(n9437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__14255.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__14256 (.I0(n9355), .I1(n9436), .I2(n9437), .I3(\i2c_config_index[6] ), 
            .O(n9438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__14256.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__14257 (.I0(n9129), .I1(n9081), .I2(n9183), .I3(n9056), 
            .O(n9439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__14257.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__14258 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[5] ), .O(n9440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he33f */ ;
    defparam LUT__14258.LUTMASK = 16'he33f;
    EFX_LUT4 LUT__14259 (.I0(n9440), .I1(\i2c_config_index[4] ), .I2(n9197), 
            .I3(\i2c_config_index[3] ), .O(n9441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__14259.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__14260 (.I0(n9441), .I1(n9439), .I2(n9261), .I3(n9143), 
            .O(n9442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__14260.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__14261 (.I0(n9438), .I1(n9442), .I2(n9434), .I3(n9044), 
            .O(n9443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__14261.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__14262 (.I0(n9137), .I1(\u_i2c_timing_ctrl_16bit/i2c_wdata[5] ), 
            .I2(n9443), .I3(n9135), .O(\u_i2c_timing_ctrl_16bit/n378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__14262.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__14263 (.I0(n9104), .I1(n9094), .I2(n9072), .O(n9444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14263.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14264 (.I0(n9101), .I1(n9325), .I2(\i2c_config_index[0] ), 
            .I3(n9444), .O(n9445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__14264.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__14265 (.I0(n9129), .I1(n9174), .I2(\i2c_config_index[3] ), 
            .O(n9446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14265.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14266 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[2] ), .O(n9447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1700 */ ;
    defparam LUT__14266.LUTMASK = 16'h1700;
    EFX_LUT4 LUT__14267 (.I0(n9446), .I1(n9447), .I2(n9445), .I3(\i2c_config_index[5] ), 
            .O(n9448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__14267.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__14268 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[2] ), .I3(n9196), .O(n9449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14268.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14269 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[5] ), .O(n9450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haf74 */ ;
    defparam LUT__14269.LUTMASK = 16'haf74;
    EFX_LUT4 LUT__14270 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[5] ), 
            .I2(\i2c_config_index[4] ), .I3(n9192), .O(n9451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00 */ ;
    defparam LUT__14270.LUTMASK = 16'h2c00;
    EFX_LUT4 LUT__14271 (.I0(n9450), .I1(n9066), .I2(n9451), .I3(n9017), 
            .O(n9452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14271.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14272 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n9453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ea3 */ ;
    defparam LUT__14272.LUTMASK = 16'h3ea3;
    EFX_LUT4 LUT__14273 (.I0(n9453), .I1(n9217), .I2(n9202), .I3(\i2c_config_index[7] ), 
            .O(n9454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__14273.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__14274 (.I0(n9454), .I1(\i2c_config_index[6] ), .I2(n9449), 
            .I3(n9452), .O(n9455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__14274.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__14275 (.I0(n9063), .I1(n9448), .I2(n9092), .I3(n9455), 
            .O(n9456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__14275.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__14276 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[3] ), .O(n9457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h83fa */ ;
    defparam LUT__14276.LUTMASK = 16'h83fa;
    EFX_LUT4 LUT__14277 (.I0(n9282), .I1(n9254), .I2(n9129), .I3(n9258), 
            .O(n9458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14277.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14278 (.I0(\i2c_config_index[1] ), .I1(n9457), .I2(n9458), 
            .O(n9459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__14278.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__14279 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[3] ), .O(n9460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfed3 */ ;
    defparam LUT__14279.LUTMASK = 16'hfed3;
    EFX_LUT4 LUT__14280 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[0] ), .O(n9461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdfe */ ;
    defparam LUT__14280.LUTMASK = 16'hbdfe;
    EFX_LUT4 LUT__14281 (.I0(n9461), .I1(n9460), .I2(\i2c_config_index[4] ), 
            .O(n9462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14281.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14282 (.I0(n9462), .I1(n9459), .I2(\i2c_config_index[5] ), 
            .I3(n9261), .O(n9463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__14282.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__14283 (.I0(n9214), .I1(n9067), .I2(n9083), .I3(n9019), 
            .O(n9464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e00 */ ;
    defparam LUT__14283.LUTMASK = 16'h3e00;
    EFX_LUT4 LUT__14284 (.I0(n9464), .I1(n9405), .I2(n9409), .O(n9465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14284.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14285 (.I0(n9279), .I1(n9019), .I2(n9017), .O(n9466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14285.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14286 (.I0(n9466), .I1(n9465), .I2(n9044), .I3(n9046), 
            .O(n9467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf530 */ ;
    defparam LUT__14286.LUTMASK = 16'hf530;
    EFX_LUT4 LUT__14287 (.I0(n9463), .I1(n9456), .I2(n9467), .O(n9468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__14287.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__14288 (.I0(n9137), .I1(\u_i2c_timing_ctrl_16bit/i2c_wdata[6] ), 
            .I2(n9468), .I3(n9135), .O(\u_i2c_timing_ctrl_16bit/n377 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f44 */ ;
    defparam LUT__14288.LUTMASK = 16'h0f44;
    EFX_LUT4 LUT__14289 (.I0(n9255), .I1(n9087), .I2(\i2c_config_index[4] ), 
            .O(n9469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14289.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14290 (.I0(n9113), .I1(n9052), .I2(\i2c_config_index[3] ), 
            .O(n9470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3 */ ;
    defparam LUT__14290.LUTMASK = 16'he3e3;
    EFX_LUT4 LUT__14291 (.I0(n9470), .I1(n9118), .I2(\i2c_config_index[5] ), 
            .O(n9471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14291.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14292 (.I0(n9182), .I1(n9469), .I2(n9471), .O(n9472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__14292.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__14293 (.I0(n9108), .I1(n9019), .I2(n9472), .I3(\i2c_config_index[7] ), 
            .O(n9473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077 */ ;
    defparam LUT__14293.LUTMASK = 16'hf077;
    EFX_LUT4 LUT__14294 (.I0(n9202), .I1(n9473), .I2(n9044), .I3(\i2c_config_index[6] ), 
            .O(n9474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__14294.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__14295 (.I0(\i2c_config_index[7] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[2] ), .O(n9475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe15 */ ;
    defparam LUT__14295.LUTMASK = 16'hfe15;
    EFX_LUT4 LUT__14296 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[5] ), .O(n9476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbffd */ ;
    defparam LUT__14296.LUTMASK = 16'hbffd;
    EFX_LUT4 LUT__14297 (.I0(n9476), .I1(n9217), .I2(n9475), .I3(\i2c_config_index[7] ), 
            .O(n9477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__14297.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__14298 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n9478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7fe */ ;
    defparam LUT__14298.LUTMASK = 16'he7fe;
    EFX_LUT4 LUT__14299 (.I0(n9478), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[5] ), 
            .O(n9479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14299.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14300 (.I0(\i2c_config_index[0] ), .I1(n9479), .I2(n9477), 
            .I3(\i2c_config_index[7] ), .O(n9480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f31 */ ;
    defparam LUT__14300.LUTMASK = 16'h0f31;
    EFX_LUT4 LUT__14301 (.I0(n9190), .I1(n9069), .I2(n9234), .O(n9481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14301.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14302 (.I0(n9234), .I1(n9053), .I2(\i2c_config_index[3] ), 
            .I3(\i2c_config_index[5] ), .O(n9482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haff3 */ ;
    defparam LUT__14302.LUTMASK = 16'haff3;
    EFX_LUT4 LUT__14303 (.I0(n9254), .I1(n9282), .I2(n9481), .I3(n9482), 
            .O(n9483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__14303.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__14304 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[5] ), .I3(n9254), .O(n9484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b00 */ ;
    defparam LUT__14304.LUTMASK = 16'h2b00;
    EFX_LUT4 LUT__14305 (.I0(n9484), .I1(n9483), .I2(\i2c_config_index[4] ), 
            .O(n9485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__14305.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__14306 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[1] ), .O(n9486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb70d */ ;
    defparam LUT__14306.LUTMASK = 16'hb70d;
    EFX_LUT4 LUT__14307 (.I0(\i2c_config_index[3] ), .I1(n9053), .I2(n9486), 
            .I3(n9098), .O(n9487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__14307.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__14308 (.I0(n9487), .I1(n9485), .I2(\i2c_config_index[7] ), 
            .I3(n9480), .O(n9488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__14308.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__14309 (.I0(\i2c_config_index[6] ), .I1(n9488), .I2(\i2c_config_index[7] ), 
            .I3(n9044), .O(n9489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__14309.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__14310 (.I0(n9474), .I1(n9489), .I2(n9046), .O(n9490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14310.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14311 (.I0(n9137), .I1(n9490), .I2(n9135), .I3(\u_i2c_timing_ctrl_16bit/i2c_wdata[7] ), 
            .O(\u_i2c_timing_ctrl_16bit/n376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcdc0 */ ;
    defparam LUT__14311.LUTMASK = 16'hcdc0;
    EFX_LUT4 LUT__14312 (.I0(n4508), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[2] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14312.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14313 (.I0(n4506), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[3] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14313.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14314 (.I0(n4504), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[4] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14314.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14315 (.I0(n4502), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[5] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14315.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14316 (.I0(n4500), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[6] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14316.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14317 (.I0(n4498), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[7] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14317.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14318 (.I0(n4496), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[8] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14318.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14319 (.I0(n4494), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[9] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14319.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14320 (.I0(n4492), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[10] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14320.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14321 (.I0(n4490), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[11] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14321.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14322 (.I0(n4488), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[12] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14322.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14323 (.I0(n4486), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[13] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14323.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14324 (.I0(n4484), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[14] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14324.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14325 (.I0(n4482), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[15] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14325.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14326 (.I0(n4480), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[16] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14326.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14327 (.I0(n4478), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[17] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14327.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14328 (.I0(n4476), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[18] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14328.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14329 (.I0(n4474), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[19] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14329.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14330 (.I0(n4472), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[20] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14330.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14331 (.I0(n4470), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[21] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14331.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14332 (.I0(n4468), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[22] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14332.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14333 (.I0(n4466), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[23] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14333.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14334 (.I0(n4464), .I1(\u_i2c_timing_ctrl_16bit/delay_cnt[24] ), 
            .I2(n9152), .O(\u_i2c_timing_ctrl_16bit/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14334.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14335 (.I0(\u_i2c_timing_ctrl_16bit/delay_cnt[25] ), .I1(n9151), 
            .I2(\u_i2c_timing_ctrl_16bit/delay_cnt[26] ), .I3(n4462), .O(\u_i2c_timing_ctrl_16bit/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfa0 */ ;
    defparam LUT__14335.LUTMASK = 16'hbfa0;
    EFX_LUT4 LUT__14336 (.I0(n9152), .I1(n4461), .O(\u_i2c_timing_ctrl_16bit/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__14336.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__14337 (.I0(n4383), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[11] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14337.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14338 (.I0(n4384), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[10] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14338.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14339 (.I0(n4386), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[9] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14339.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14340 (.I0(cmos_href), .I1(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .I2(\u_Sensor_Image_XYCrop_0/image_ypos[0] ), .O(\u_Sensor_Image_XYCrop_0/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__14340.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__14341 (.I0(n4388), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[8] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n45 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14341.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14342 (.I0(n4390), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[7] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14342.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14343 (.I0(n4392), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[6] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14343.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14344 (.I0(n4394), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[5] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14344.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14345 (.I0(n4396), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[4] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14345.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14346 (.I0(n4398), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[3] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14346.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14347 (.I0(n4400), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[2] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14347.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14348 (.I0(\u_Sensor_Image_XYCrop_0/image_ypos[4] ), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[5] ), 
            .I2(\u_Sensor_Image_XYCrop_0/image_ypos[7] ), .I3(\u_Sensor_Image_XYCrop_0/image_ypos[6] ), 
            .O(n9491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__14348.LUTMASK = 16'he000;
    EFX_LUT4 LUT__14349 (.I0(\u_Sensor_Image_XYCrop_0/image_xpos[10] ), .I1(\u_Sensor_Image_XYCrop_0/image_xpos[9] ), 
            .I2(\u_Sensor_Image_XYCrop_0/image_xpos[11] ), .O(n9492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__14349.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__14350 (.I0(n9492), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[11] ), 
            .I2(\u_Sensor_Image_XYCrop_0/image_ypos[10] ), .I3(cmos_href), 
            .O(n9493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14350.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14351 (.I0(n9491), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[8] ), 
            .I2(\u_Sensor_Image_XYCrop_0/image_ypos[9] ), .I3(n9493), .O(\u_Sensor_Image_XYCrop_0/w_image_out_href )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__14351.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__14352 (.I0(n541), .I1(\u_Sensor_Image_XYCrop_0/image_ypos[1] ), 
            .I2(cmos_href), .I3(\u_Sensor_Image_XYCrop_0/image_in_href_r ), 
            .O(\u_Sensor_Image_XYCrop_0/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14352.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14353 (.I0(DdrCtrl_ARVALID_0), .I1(DdrCtrl_AWVALID_0), 
            .I2(DdrCtrl_ATYPE_0), .O(n9494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14353.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14354 (.I0(n9494), .I1(DdrCtrl_AREADY_0), .I2(\axi4_awar_mux/rs_req[1] ), 
            .I3(\axi4_awar_mux/rs_req[0] ), .O(\axi4_awar_mux/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__14354.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__14355 (.I0(\axi4_awar_mux/rs_req[1] ), .I1(\axi4_awar_mux/rs_req[0] ), 
            .I2(DdrCtrl_AREADY_0), .O(\axi4_awar_mux/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14355.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14356 (.I0(\axi4_awar_mux/rs_req[0] ), .I1(\axi4_awar_mux/rs_req[1] ), 
            .I2(n9494), .O(n9495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14356.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14357 (.I0(\axi4_awar_mux/n131 ), .I1(DdrCtrl_AVALID_0), 
            .I2(n9495), .O(\axi4_awar_mux/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__14357.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__14358 (.I0(\axi4_awar_mux/rs_req[0] ), .I1(\axi4_awar_mux/rs_req[1] ), 
            .I2(DdrCtrl_ATYPE_0), .O(\axi4_awar_mux/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__14358.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__14359 (.I0(n9494), .I1(DdrCtrl_AREADY_0), .I2(\axi4_awar_mux/rs_req[1] ), 
            .I3(\axi4_awar_mux/rs_req[0] ), .O(\axi4_awar_mux/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__14359.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__14360 (.I0(\DdrCtrl_AWADDR_0[23] ), .I1(\u_axi4_ctrl_0/r_wframe_index_last[1] ), 
            .I2(\u_axi4_ctrl_0/r_rframe_inc ), .I3(\u_axi4_ctrl_0/r_wframe_inc ), 
            .O(\u_axi4_ctrl_0/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14360.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14361 (.I0(\DdrCtrl_AWADDR_0[23] ), .I1(\u_axi4_ctrl_0/r_wframe_index_last[1] ), 
            .I2(\u_axi4_ctrl_0/r_wframe_inc ), .O(n9496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14361.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14362 (.I0(\DdrCtrl_ARADDR_0[23] ), .I1(n9496), .I2(\u_axi4_ctrl_0/r_rframe_inc ), 
            .O(\u_axi4_ctrl_0/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__14362.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__14363 (.I0(\DdrCtrl_AWADDR_0[22] ), .I1(\u_axi4_ctrl_0/r_wframe_index_last[0] ), 
            .I2(\u_axi4_ctrl_0/r_wframe_inc ), .O(n9497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14363.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14364 (.I0(\DdrCtrl_ARADDR_0[22] ), .I1(n9497), .I2(\u_axi4_ctrl_0/r_rframe_inc ), 
            .O(\u_axi4_ctrl_0/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__14364.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__14365 (.I0(\DdrCtrl_AWADDR_0[22] ), .I1(\u_axi4_ctrl_0/r_wframe_index_last[0] ), 
            .I2(\u_axi4_ctrl_0/r_rframe_inc ), .I3(\u_axi4_ctrl_0/r_wframe_inc ), 
            .O(\u_axi4_ctrl_0/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__14365.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__14366 (.I0(n4283), .I1(n4284), .I2(n4286), .I3(n4288), 
            .O(n9498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14366.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14367 (.I0(n4290), .I1(n9498), .O(n9499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14367.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14369 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .O(n9501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14369.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14371 (.I0(\u_axi4_ctrl_0/rs_w[1] ), .I1(DdrCtrl_WREADY_0), 
            .I2(DdrCtrl_WLAST_0), .O(n9503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14371.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14372 (.I0(\u_axi4_ctrl_0/rc_w_eof[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9503), .I3(\u_axi4_ctrl_0/rs_w[0] ), .O(n9504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__14372.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__14373 (.I0(\u_axi4_ctrl_0/r_weof_pending ), .I1(n9499), 
            .I2(n9501), .I3(n9504), .O(\u_axi4_ctrl_0/n265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__14373.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__14374 (.I0(n4304), .I1(n4306), .I2(n4308), .I3(n4310), 
            .O(n9505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14374.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14375 (.I0(n4296), .I1(n4298), .I2(n4300), .I3(n4302), 
            .O(n9506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14375.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14376 (.I0(n961), .I1(n4295), .I2(n9505), .I3(n9506), 
            .O(n9507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14376.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14377 (.I0(DdrCtrl_WREADY_0), .I1(DdrCtrl_WVALID_0), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .I3(n9507), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__14377.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__14378 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I3(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .O(n9508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0990 */ ;
    defparam LUT__14378.LUTMASK = 16'h0990;
    EFX_LUT4 LUT__14379 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .I2(n9508), .O(n9509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__14379.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__14380 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] ), 
            .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] ), .I3(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .O(n9510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14380.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14381 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] ), .I3(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .O(n9511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14381.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14382 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] ), 
            .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] ), .I3(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .O(n9512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14382.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14383 (.I0(n9509), .I1(n9510), .I2(n9511), .I3(n9512), 
            .O(n9513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14383.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14384 (.I0(r_XYCrop0_frame_href), .I1(r_XYCrop0_frame_de), 
            .O(n9514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14384.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14385 (.I0(n9514), .I1(\u_axi4_ctrl_0/rc_wfifo_we[0] ), 
            .I2(\u_axi4_ctrl_0/rc_wfifo_we[1] ), .O(n9515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14385.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14386 (.I0(n9513), .I1(n9515), .I2(\u_axi4_ctrl_0/rc_wfifo_we[2] ), 
            .I3(\u_axi4_ctrl_0/rc_wfifo_we[3] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__14386.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__14387 (.I0(\u_axi4_ctrl_0/rs_w[1] ), .I1(\u_axi4_ctrl_0/rs_w[0] ), 
            .O(n9516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14387.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14388 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[0] ), .O(\u_axi4_ctrl_0/n290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14388.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14389 (.I0(\u_axi4_ctrl_0/rc_w_eof[0] ), .I1(n9516), .O(\u_axi4_ctrl_0/n291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14389.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14390 (.I0(\u_axi4_ctrl_0/w_wfifo_empty ), .I1(\u_axi4_ctrl_0/r_weof_pending ), 
            .I2(n9499), .I3(n9501), .O(n9517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__14390.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__14391 (.I0(DdrCtrl_AWREADY_0), .I1(DdrCtrl_AWVALID_0), 
            .I2(n9517), .O(\u_axi4_ctrl_0/n258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__14391.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__14392 (.I0(n9503), .I1(\u_axi4_ctrl_0/rs_w[0] ), .O(n9518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14392.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14393 (.I0(DdrCtrl_WVALID_0), .I1(n9517), .I2(n9518), 
            .O(\u_axi4_ctrl_0/n260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__14393.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__14394 (.I0(\u_axi4_ctrl_0/rs_w[1] ), .I1(\Axi0ResetReg[2] ), 
            .O(n9519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14394.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14395 (.I0(n546), .I1(\u_axi4_ctrl_0/rs_w[0] ), .I2(\u_axi4_ctrl_0/rc_burst[0] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14395.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14396 (.I0(\u_axi4_ctrl_0/r_wframe_sync[0] ), .I1(\u_axi4_ctrl_0/r_wframe_sync[1] ), 
            .I2(\u_axi4_ctrl_0/r_weof_pending ), .I3(n9516), .O(\u_axi4_ctrl_0/n267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__14396.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__14397 (.I0(n9501), .I1(n9499), .I2(\u_axi4_ctrl_0/r_weof_pending ), 
            .I3(\u_axi4_ctrl_0/w_wfifo_empty ), .O(\u_axi4_ctrl_0/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14397.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14399 (.I0(n9514), .I1(\u_axi4_ctrl_0/rc_wfifo_we[0] ), 
            .O(\u_axi4_ctrl_0/n2649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14399.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14400 (.I0(\u_axi4_ctrl_0/rfifo_cnt[1] ), .I1(\u_axi4_ctrl_0/rfifo_cnt[0] ), 
            .I2(\u_axi4_ctrl_0/rfifo_cnt[2] ), .I3(\u_axi4_ctrl_0/rfifo_cnt[3] ), 
            .O(n9520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14400.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14401 (.I0(\u_axi4_ctrl_0/rfifo_cnt[4] ), .I1(n9520), 
            .O(\u_axi4_ctrl_0/equal_138/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14401.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14402 (.I0(\u_axi4_ctrl_0/equal_138/n9 ), .I1(n4281), 
            .O(\u_axi4_ctrl_0/n1074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14402.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14403 (.I0(lcd_vs), .I1(\u_axi4_ctrl_0/rframe_vsync_dly ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl_0/n2551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__14403.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__14404 (.I0(\u_axi4_ctrl_0/equal_138/n9 ), .I1(n978), .O(\u_axi4_ctrl_0/n1075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14404.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14405 (.I0(\u_axi4_ctrl_0/rfifo_rst ), .I1(\Axi0ResetReg[2] ), 
            .O(\u_axi4_ctrl_0/w_rfifo_rst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14405.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14406 (.I0(\u_axi4_ctrl_0/rc_rfifo_rd[0] ), .I1(lcd_request), 
            .O(\u_axi4_ctrl_0/n2670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14406.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14409 (.I0(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[1] ), .I1(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[0] ), 
            .O(\u_axi4_ctrl_0/equal_160/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14409.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14412 (.I0(\DdrCtrl_ARADDR_0[13] ), .I1(\DdrCtrl_ARADDR_0[14] ), 
            .I2(\DdrCtrl_ARADDR_0[15] ), .I3(\DdrCtrl_ARADDR_0[16] ), .O(n9523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14412.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14413 (.I0(\DdrCtrl_ARADDR_0[18] ), .I1(\DdrCtrl_ARADDR_0[19] ), 
            .I2(\DdrCtrl_ARADDR_0[20] ), .O(n9524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14413.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14414 (.I0(\DdrCtrl_ARADDR_0[21] ), .I1(n4220), .I2(n4221), 
            .I3(\u_axi4_ctrl_0/rfifo_wr_rst_busy_dly[15] ), .O(n9525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14414.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14415 (.I0(\DdrCtrl_ARADDR_0[17] ), .I1(n9523), .I2(n9524), 
            .I3(n9525), .O(n9526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__14415.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__14416 (.I0(DdrCtrl_ARVALID_0), .I1(\u_axi4_ctrl_0/r_rd_pend ), 
            .O(n9527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14416.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14417 (.I0(n9527), .I1(n9526), .I2(\u_axi4_ctrl_0/rd_state.S_READ_IDLE ), 
            .I3(\u_axi4_ctrl_0/rd_state.S_READ_DATA ), .O(n9528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf5cf */ ;
    defparam LUT__14417.LUTMASK = 16'hf5cf;
    EFX_LUT4 LUT__14418 (.I0(n9528), .I1(\u_axi4_ctrl_0/rd_state.S_READ_ADDR ), 
            .O(\u_axi4_ctrl_0/n1730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14418.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14419 (.I0(\u_axi4_ctrl_0/rd_state.S_READ_ADDR ), .I1(\u_axi4_ctrl_0/rd_state.S_READ_DATA ), 
            .I2(n9526), .I3(\u_axi4_ctrl_0/rd_state.S_READ_IDLE ), .O(\u_axi4_ctrl_0/select_190/Select_1/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14419.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14420 (.I0(\u_axi4_ctrl_0/rd_state.S_READ_IDLE ), .I1(\u_axi4_ctrl_0/rd_state.S_READ_ADDR ), 
            .I2(\u_axi4_ctrl_0/rd_state.S_READ_DATA ), .O(\u_axi4_ctrl_0/equal_189/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__14420.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__14421 (.I0(\u_axi4_ctrl_0/rd_state.S_READ_IDLE ), .I1(\u_axi4_ctrl_0/rd_state.S_READ_DATA ), 
            .I2(\u_axi4_ctrl_0/rd_state.S_READ_ADDR ), .O(n9529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14421.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14422 (.I0(n9527), .I1(\u_axi4_ctrl_0/equal_189/n5 ), 
            .I2(n9529), .O(\u_axi4_ctrl_0/n1732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf1f1 */ ;
    defparam LUT__14422.LUTMASK = 16'hf1f1;
    EFX_LUT4 LUT__14423 (.I0(DdrCtrl_ARREADY_0), .I1(DdrCtrl_ARVALID_0), 
            .I2(n9529), .O(\u_axi4_ctrl_0/n1733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__14423.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__14424 (.I0(DdrCtrl_RLAST_0), .I1(DdrCtrl_RVALID_0), .I2(\u_axi4_ctrl_0/r_rd_pend ), 
            .I3(n9529), .O(\u_axi4_ctrl_0/n1734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__14424.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__14431 (.I0(\u_axi4_ctrl_0/rc_w_eof[0] ), .I1(\u_axi4_ctrl_0/rs_w[0] ), 
            .O(n9530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14431.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14432 (.I0(\u_axi4_ctrl_0/rs_w[1] ), .I1(n9530), .I2(n9518), 
            .I3(\u_axi4_ctrl_0/n266 ), .O(\u_axi4_ctrl_0/n264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2 */ ;
    defparam LUT__14432.LUTMASK = 16'hfff2;
    EFX_LUT4 LUT__14433 (.I0(\DdrCtrl_ARADDR_0[23] ), .I1(\DdrCtrl_AWADDR_0[23] ), 
            .O(n9531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14433.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14434 (.I0(n9531), .I1(\DdrCtrl_ARADDR_0[22] ), .I2(\u_axi4_ctrl_0/r_wframe_inc ), 
            .I3(\DdrCtrl_AWADDR_0[22] ), .O(\u_axi4_ctrl_0/n2777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2fb0 */ ;
    defparam LUT__14434.LUTMASK = 16'h2fb0;
    EFX_LUT4 LUT__14435 (.I0(n9501), .I1(\u_axi4_ctrl_0/r_w_rst ), .I2(\u_axi4_ctrl_0/n266 ), 
            .O(\u_axi4_ctrl_0/n256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf1f1 */ ;
    defparam LUT__14435.LUTMASK = 16'hf1f1;
    EFX_LUT4 LUT__14436 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[1] ), .O(\u_axi4_ctrl_0/n289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14436.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14437 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[2] ), .O(\u_axi4_ctrl_0/n288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14437.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14438 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[3] ), .O(\u_axi4_ctrl_0/n287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14438.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14439 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[4] ), .O(\u_axi4_ctrl_0/n286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14439.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14440 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[5] ), .O(\u_axi4_ctrl_0/n285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14440.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14441 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[6] ), .O(\u_axi4_ctrl_0/n284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14441.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14442 (.I0(n9516), .I1(\DdrCtrl_AWADDR_0[7] ), .O(\u_axi4_ctrl_0/n283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14442.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14443 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\DdrCtrl_AWADDR_0[8] ), 
            .I2(\u_axi4_ctrl_0/rs_w[1] ), .O(\u_axi4_ctrl_0/n282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1c1c */ ;
    defparam LUT__14443.LUTMASK = 16'h1c1c;
    EFX_LUT4 LUT__14444 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(\DdrCtrl_AWADDR_0[8] ), .I3(\DdrCtrl_AWADDR_0[9] ), .O(\u_axi4_ctrl_0/n281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14444.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14445 (.I0(\DdrCtrl_AWADDR_0[8] ), .I1(\DdrCtrl_AWADDR_0[9] ), 
            .O(n9532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14445.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14446 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9532), .I3(\DdrCtrl_AWADDR_0[10] ), .O(\u_axi4_ctrl_0/n280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14446.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14447 (.I0(\u_axi4_ctrl_0/rs_w[1] ), .I1(n9532), .I2(\DdrCtrl_AWADDR_0[10] ), 
            .O(n9533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14447.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14448 (.I0(n9516), .I1(n9533), .I2(\DdrCtrl_AWADDR_0[11] ), 
            .O(\u_axi4_ctrl_0/n279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__14448.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__14449 (.I0(n9532), .I1(\DdrCtrl_AWADDR_0[10] ), .I2(\DdrCtrl_AWADDR_0[11] ), 
            .O(n9534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14449.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14450 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9534), .I3(\DdrCtrl_AWADDR_0[12] ), .O(\u_axi4_ctrl_0/n278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14450.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14451 (.I0(n9534), .I1(\DdrCtrl_AWADDR_0[12] ), .O(n9535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14451.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14452 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9535), .I3(\DdrCtrl_AWADDR_0[13] ), .O(\u_axi4_ctrl_0/n277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14452.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14453 (.I0(n9535), .I1(\DdrCtrl_AWADDR_0[13] ), .O(n9536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14453.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14454 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9536), .I3(\DdrCtrl_AWADDR_0[14] ), .O(\u_axi4_ctrl_0/n276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14454.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14455 (.I0(n9536), .I1(\DdrCtrl_AWADDR_0[14] ), .O(n9537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14455.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14456 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9537), .I3(\DdrCtrl_AWADDR_0[15] ), .O(\u_axi4_ctrl_0/n275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14456.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14457 (.I0(n9537), .I1(\DdrCtrl_AWADDR_0[15] ), .O(n9538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14457.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14458 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9538), .I3(\DdrCtrl_AWADDR_0[16] ), .O(\u_axi4_ctrl_0/n274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14458.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14459 (.I0(n9538), .I1(\DdrCtrl_AWADDR_0[16] ), .O(n9539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14459.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14460 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9539), .I3(\DdrCtrl_AWADDR_0[17] ), .O(\u_axi4_ctrl_0/n273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14460.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14461 (.I0(n9539), .I1(\DdrCtrl_AWADDR_0[17] ), .O(n9540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14461.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14462 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9540), .I3(\DdrCtrl_AWADDR_0[18] ), .O(\u_axi4_ctrl_0/n272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14462.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14463 (.I0(n9540), .I1(\DdrCtrl_AWADDR_0[18] ), .O(n9541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14463.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14464 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9541), .I3(\DdrCtrl_AWADDR_0[19] ), .O(\u_axi4_ctrl_0/n271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14464.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14465 (.I0(n9541), .I1(\DdrCtrl_AWADDR_0[19] ), .O(n9542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14465.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14466 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9542), .I3(\DdrCtrl_AWADDR_0[20] ), .O(\u_axi4_ctrl_0/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14466.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14467 (.I0(n9542), .I1(\DdrCtrl_AWADDR_0[20] ), .O(n9543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14467.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14468 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(\u_axi4_ctrl_0/rs_w[1] ), 
            .I2(n9543), .I3(\DdrCtrl_AWADDR_0[21] ), .O(\u_axi4_ctrl_0/n269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3740 */ ;
    defparam LUT__14468.LUTMASK = 16'h3740;
    EFX_LUT4 LUT__14469 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(n4381), .I2(\u_axi4_ctrl_0/rc_burst[1] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n345 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14469.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14470 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(n4379), .I2(\u_axi4_ctrl_0/rc_burst[2] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14470.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14471 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(n4377), .I2(\u_axi4_ctrl_0/rc_burst[3] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14471.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14472 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(n4375), .I2(\u_axi4_ctrl_0/rc_burst[4] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14472.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14473 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(n4373), .I2(\u_axi4_ctrl_0/rc_burst[5] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14473.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14474 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(n4371), .I2(\u_axi4_ctrl_0/rc_burst[6] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14474.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14475 (.I0(\u_axi4_ctrl_0/rs_w[0] ), .I1(n4370), .I2(\u_axi4_ctrl_0/rc_burst[7] ), 
            .I3(n9519), .O(\u_axi4_ctrl_0/n339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__14475.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__14483 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[8] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[16] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14483.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14484 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[9] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[17] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14484.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14485 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[10] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[18] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14485.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14486 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[11] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[19] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14486.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14487 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[12] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[20] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14487.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14488 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[13] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[21] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14488.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14489 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[14] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[22] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14489.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14490 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[15] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[23] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14490.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14491 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[16] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[24] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14491.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14492 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[17] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[25] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14492.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14493 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[18] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[26] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14493.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14494 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[19] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[27] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14494.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14495 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[20] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[28] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14495.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14496 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[21] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[29] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14496.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14497 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[22] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[30] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14497.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14498 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[23] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[31] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14498.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14499 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[24] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[32] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14499.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14500 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[25] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[33] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14500.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14501 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[26] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[34] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14501.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14502 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[27] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[35] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14502.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14503 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[28] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[36] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14503.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14504 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[29] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[37] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14504.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14505 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[30] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[38] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14505.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14506 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[31] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[39] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14506.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14507 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[32] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[40] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14507.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14508 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[33] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[41] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14508.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14509 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[34] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[42] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14509.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14510 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[35] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[43] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14510.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14511 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[36] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[44] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14511.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14512 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[37] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[45] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14512.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14513 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[38] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[46] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14513.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14514 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[39] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[47] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14514.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14515 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[40] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[48] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14515.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14516 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[41] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[49] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14516.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14517 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[42] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[50] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14517.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14518 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[43] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[51] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14518.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14519 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[44] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[52] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14519.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14520 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[45] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[53] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n729 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14520.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14521 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[46] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[54] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14521.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14522 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[47] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[55] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n727 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14522.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14523 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[48] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[56] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14523.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14524 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[49] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[57] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14524.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14525 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[50] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[58] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n724 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14525.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14526 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[51] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[59] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n723 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14526.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14527 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[52] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[60] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14527.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14528 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[53] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[61] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n721 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14528.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14529 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[54] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[62] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14529.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14530 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[55] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[63] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n719 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14530.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14531 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[56] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[64] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14531.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14532 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[57] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[65] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n717 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14532.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14533 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[58] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[66] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14533.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14534 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[59] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[67] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14534.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14535 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[60] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[68] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14535.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14536 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[61] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[69] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14536.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14537 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[62] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[70] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14537.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14538 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[63] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[71] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14538.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14539 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[64] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[72] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14539.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14540 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[65] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[73] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n709 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14540.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14541 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[66] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[74] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14541.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14542 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[67] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[75] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n707 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14542.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14543 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[68] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[76] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n706 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14543.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14544 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[69] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[77] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14544.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14545 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[70] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[78] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14545.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14546 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[71] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[79] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14546.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14547 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[72] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[80] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14547.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14548 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[73] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[81] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n701 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14548.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14549 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[74] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[82] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14549.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14550 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[75] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[83] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14550.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14551 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[76] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[84] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14551.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14552 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[77] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[85] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14552.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14553 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[78] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[86] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14553.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14554 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[79] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[87] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14554.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14555 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[80] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[88] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14555.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14556 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[81] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[89] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14556.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14557 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[82] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[90] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14557.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14558 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[83] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[91] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14558.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14559 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[84] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[92] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14559.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14560 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[85] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[93] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14560.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14561 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[86] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[94] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14561.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14562 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[87] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[95] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14562.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14563 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[88] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[96] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14563.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14564 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[89] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[97] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14564.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14565 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[90] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[98] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14565.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14566 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[91] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[99] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14566.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14567 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[92] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[100] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14567.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14568 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[93] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[101] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14568.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14569 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[94] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[102] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14569.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14570 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[95] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[103] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n679 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14570.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14571 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[96] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[104] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14571.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14572 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[97] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[105] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14572.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14573 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[98] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[106] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n676 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14573.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14574 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[99] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[107] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n675 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14574.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14575 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[100] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[108] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n674 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14575.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14576 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[101] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[109] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14576.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14577 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[102] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[110] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14577.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14578 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[103] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[111] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n671 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14578.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14579 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[104] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[112] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14579.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14580 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[105] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[113] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n669 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14580.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14581 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[106] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[114] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n668 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14581.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14582 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[107] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[115] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14582.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14583 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[108] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[116] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14583.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14584 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[109] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[117] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14584.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14585 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[110] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[118] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n664 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14585.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14586 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[111] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[119] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14586.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14587 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[112] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[120] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n662 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14587.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14588 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[113] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[121] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14588.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14589 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[114] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[122] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14589.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14590 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[115] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[123] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14590.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14591 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[116] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[124] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14591.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14592 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[117] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[125] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n657 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14592.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14593 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[118] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[126] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14593.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14594 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[119] ), .I1(\u_axi4_ctrl_0/r_wfifo_wdata[127] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n655 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14594.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14595 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[120] ), .I1(\r_XYCrop0_frame_Gray[0] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n654 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14595.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14596 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[121] ), .I1(\r_XYCrop0_frame_Gray[1] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n653 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14596.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14597 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[122] ), .I1(\r_XYCrop0_frame_Gray[2] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14597.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14598 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[123] ), .I1(\r_XYCrop0_frame_Gray[3] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n651 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14598.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14599 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[124] ), .I1(\r_XYCrop0_frame_Gray[4] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n650 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14599.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14600 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[125] ), .I1(\r_XYCrop0_frame_Gray[5] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14600.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14601 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[126] ), .I1(\r_XYCrop0_frame_Gray[6] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14601.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14602 (.I0(\u_axi4_ctrl_0/r_wfifo_wdata[127] ), .I1(\r_XYCrop0_frame_Gray[7] ), 
            .I2(n9514), .O(\u_axi4_ctrl_0/n647 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14602.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14603 (.I0(n9514), .I1(\u_axi4_ctrl_0/rc_wfifo_we[0] ), 
            .I2(\u_axi4_ctrl_0/rc_wfifo_we[1] ), .O(\u_axi4_ctrl_0/n2656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14603.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14604 (.I0(n9515), .I1(\u_axi4_ctrl_0/rc_wfifo_we[2] ), 
            .O(\u_axi4_ctrl_0/n2661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14604.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14605 (.I0(n9515), .I1(\u_axi4_ctrl_0/rc_wfifo_we[2] ), 
            .I2(\u_axi4_ctrl_0/rc_wfifo_we[3] ), .O(\u_axi4_ctrl_0/n2666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14605.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14606 (.I0(\u_axi4_ctrl_0/rc_rfifo_rd[0] ), .I1(\u_axi4_ctrl_0/rc_rfifo_rd[1] ), 
            .I2(\u_axi4_ctrl_0/rc_rfifo_rd[2] ), .I3(lcd_request), .O(n9544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14606.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14607 (.I0(n4244), .I1(n4246), .I2(n4248), .I3(n4250), 
            .O(n9545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14607.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14608 (.I0(n4236), .I1(n4238), .I2(n4240), .I3(n4242), 
            .O(n9546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14608.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14609 (.I0(n1208), .I1(n4235), .I2(n9545), .I3(n9546), 
            .O(n9547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14609.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14610 (.I0(\u_axi4_ctrl_0/w_rfifo_empty ), .I1(n9544), 
            .I2(n9547), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__14610.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__14611 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I3(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .O(n9548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0990 */ ;
    defparam LUT__14611.LUTMASK = 16'h0990;
    EFX_LUT4 LUT__14612 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] ), .I3(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .O(n9549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14612.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14613 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] ), .I3(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .O(n9550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14613.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14614 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] ), 
            .I2(n9549), .I3(n9550), .O(n9551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14614.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14615 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] ), .I3(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .O(n9552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14615.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14616 (.I0(n9551), .I1(n9552), .I2(n9548), .I3(\u_axi4_ctrl_0/rfifo_wenb ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14616.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14617 (.I0(DdrCtrl_WREADY_0), .I1(DdrCtrl_WVALID_0), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .I3(n9507), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__14617.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__14618 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14618.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14619 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14619.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14620 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14620.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14621 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14621.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14622 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14622.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14623 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14623.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14624 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14624.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14625 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14625.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14626 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14626.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14627 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14627.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14628 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14628.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14629 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14629.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14630 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14630.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14631 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14631.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14632 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14632.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14633 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14633.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14634 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14634.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14635 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14635.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14636 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14636.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14637 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n8672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14637.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14638 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[0] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n5390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14638.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14639 (.I0(n8672), .I1(n5390), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14639.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14640 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14640.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14642 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(n929), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14642.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14643 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(n954), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14643.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14644 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(n4334), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14644.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14645 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(n4332), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14645.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14646 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] ), 
            .I1(n4330), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14646.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14647 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] ), 
            .I1(n4328), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14647.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14648 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(n4326), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14648.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14649 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(n4325), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14649.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14650 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] ), 
            .I1(n958), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14650.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14651 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] ), 
            .I1(n4323), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14651.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14652 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] ), 
            .I1(n4321), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14652.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14653 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] ), 
            .I1(n4319), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14653.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14654 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] ), 
            .I1(n4317), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14654.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14655 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] ), 
            .I1(n4315), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14655.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14656 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] ), 
            .I1(n4313), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14656.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14657 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I1(n4312), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14657.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14658 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[1] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14658.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14659 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14659.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14660 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14660.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14661 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14661.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14662 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14662.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14663 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14663.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14664 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] ), .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14664.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14665 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I2(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/rd_en_int ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14665.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14666 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[2] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n8669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14666.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14667 (.I0(n8672), .I1(n8669), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14667.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14668 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[3] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n8666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14668.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14669 (.I0(n8669), .I1(n8666), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14669.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14670 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[4] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n8663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14670.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14671 (.I0(n8666), .I1(n8663), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14671.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14672 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[5] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n8660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14672.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14673 (.I0(n8663), .I1(n8660), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14673.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14674 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[6] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n8657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14674.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14675 (.I0(n8660), .I1(n8657), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14675.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14676 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/raddr[7] ), .I2(\u_axi4_ctrl_0/w_wfifo_empty ), 
            .O(n8654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14676.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14677 (.I0(n8657), .I1(n8654), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14677.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14678 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I2(\u_axi4_ctrl_0/w_wfifo_empty ), .O(n8651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14678.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14679 (.I0(n8654), .I1(n8651), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14679.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14680 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14680.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14681 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14681.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14682 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14682.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14683 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14683.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14684 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14684.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14685 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14685.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14686 (.I0(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .O(\u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14686.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14687 (.I0(\u_axi4_ctrl_0/equal_138/n9 ), .I1(n4279), 
            .O(\u_axi4_ctrl_0/n1073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14687.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14688 (.I0(\u_axi4_ctrl_0/equal_138/n9 ), .I1(n4277), 
            .O(\u_axi4_ctrl_0/n1072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14688.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14689 (.I0(\u_axi4_ctrl_0/equal_138/n9 ), .I1(n4276), 
            .O(\u_axi4_ctrl_0/n1071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14689.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14690 (.I0(\u_axi4_ctrl_0/w_rfifo_empty ), .I1(n9544), 
            .I2(n9547), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__14690.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__14691 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14691.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14692 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14692.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14693 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14693.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14694 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14694.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14695 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14695.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14696 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14696.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14697 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14697.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14698 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14698.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14699 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14699.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14700 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14700.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14701 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14701.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14702 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14702.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14703 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14703.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14704 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14704.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14705 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14705.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14706 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14706.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14707 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14707.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14708 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14708.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14709 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14709.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14710 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .O(n9553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14710.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14711 (.I0(n9553), .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[0] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] ), .I3(\u_axi4_ctrl_0/w_rfifo_empty ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__14711.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__14712 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14712.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14714 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(n1194), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14714.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14715 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(n1201), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14715.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14716 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(n4274), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14716.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14717 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(n4272), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14717.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14718 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] ), 
            .I1(n4270), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14718.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14719 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] ), 
            .I1(n4268), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14719.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14720 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(n4266), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14720.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14721 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(n4265), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/wr_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14721.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14722 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] ), 
            .I1(n1205), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14722.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14723 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] ), 
            .I1(n4263), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14723.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14724 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] ), 
            .I1(n4261), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14724.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14725 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] ), 
            .I1(n4259), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14725.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14726 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] ), 
            .I1(n4257), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14726.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14727 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] ), 
            .I1(n4255), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14727.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14728 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] ), 
            .I1(n4253), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14728.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14729 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I1(n4252), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14729.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14730 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14730.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14731 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14731.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14732 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14732.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14733 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14733.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14734 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14734.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14735 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14735.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14736 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] ), .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14736.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14737 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/rd_en_int ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/n186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14737.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14738 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .O(n9554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14738.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14739 (.I0(n9554), .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[1] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] ), .I3(\u_axi4_ctrl_0/w_rfifo_empty ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__14739.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__14740 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .O(n9555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14740.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14741 (.I0(n9555), .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[2] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] ), .I3(\u_axi4_ctrl_0/w_rfifo_empty ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__14741.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__14742 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .O(n9556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14742.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14743 (.I0(n9556), .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[3] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] ), .I3(\u_axi4_ctrl_0/w_rfifo_empty ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__14743.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__14744 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .O(n9557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14744.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14745 (.I0(n9557), .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[4] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] ), .I3(\u_axi4_ctrl_0/w_rfifo_empty ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__14745.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__14746 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .O(n9558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14746.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14747 (.I0(n9558), .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[5] ), 
            .I2(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] ), .I3(\u_axi4_ctrl_0/w_rfifo_empty ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__14747.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__14748 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[7] ), .I2(\u_axi4_ctrl_0/w_rfifo_empty ), 
            .O(n9559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__14748.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__14749 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/raddr[6] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I2(\u_axi4_ctrl_0/w_rfifo_empty ), .I3(n9559), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53 */ ;
    defparam LUT__14749.LUTMASK = 16'hac53;
    EFX_LUT4 LUT__14750 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I2(\u_axi4_ctrl_0/w_rfifo_empty ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__14750.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__14751 (.I0(n9559), .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14751.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14752 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14752.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14753 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14753.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14754 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14754.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14755 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14755.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14756 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14756.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14757 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14757.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14758 (.I0(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .O(\u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14758.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14759 (.I0(\u_axi4_ctrl_0/rc_rfifo_rd[0] ), .I1(lcd_request), 
            .I2(\u_axi4_ctrl_0/rc_rfifo_rd[1] ), .O(\u_axi4_ctrl_0/n2677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14759.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14760 (.I0(\u_axi4_ctrl_0/rc_rfifo_rd[0] ), .I1(\u_axi4_ctrl_0/rc_rfifo_rd[1] ), 
            .I2(lcd_request), .I3(\u_axi4_ctrl_0/rc_rfifo_rd[2] ), .O(\u_axi4_ctrl_0/n2682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14760.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14761 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[16] ), .I1(\lcd_data[0] ), 
            .I2(lcd_request), .O(n9560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14761.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14762 (.I0(n9560), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[0] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14762.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14763 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[17] ), .I1(\lcd_data[1] ), 
            .I2(lcd_request), .O(n9561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14763.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14764 (.I0(n9561), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[1] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14764.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14765 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[18] ), .I1(\lcd_data[2] ), 
            .I2(lcd_request), .O(n9562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14765.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14766 (.I0(n9562), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[2] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14766.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14767 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[19] ), .I1(\lcd_data[3] ), 
            .I2(lcd_request), .O(n9563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14767.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14768 (.I0(n9563), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[3] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14768.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14769 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[20] ), .I1(\lcd_data[4] ), 
            .I2(lcd_request), .O(n9564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14769.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14770 (.I0(n9564), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[4] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14770.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14771 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[21] ), .I1(\lcd_data[5] ), 
            .I2(lcd_request), .O(n9565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14771.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14772 (.I0(n9565), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[5] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14772.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14773 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[22] ), .I1(\lcd_data[6] ), 
            .I2(lcd_request), .O(n9566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14773.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14774 (.I0(n9566), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[6] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14774.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14775 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[23] ), .I1(\lcd_data[7] ), 
            .I2(lcd_request), .O(n9567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14775.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14776 (.I0(n9567), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[7] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14776.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14777 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[24] ), .I1(\lcd_data[8] ), 
            .I2(lcd_request), .O(n9568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14777.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14778 (.I0(n9568), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[8] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14778.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14779 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[25] ), .I1(\lcd_data[9] ), 
            .I2(lcd_request), .O(n9569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14779.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14780 (.I0(n9569), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[9] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14780.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14781 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[26] ), .I1(\lcd_data[10] ), 
            .I2(lcd_request), .O(n9570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14781.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14782 (.I0(n9570), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[10] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14782.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14783 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[27] ), .I1(\lcd_data[11] ), 
            .I2(lcd_request), .O(n9571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14783.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14784 (.I0(n9571), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[11] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14784.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14785 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[28] ), .I1(\lcd_data[12] ), 
            .I2(lcd_request), .O(n9572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14785.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14786 (.I0(n9572), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[12] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14786.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14787 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[29] ), .I1(\lcd_data[13] ), 
            .I2(lcd_request), .O(n9573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14787.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14788 (.I0(n9573), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[13] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14788.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14789 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[30] ), .I1(\lcd_data[14] ), 
            .I2(lcd_request), .O(n9574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14789.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14790 (.I0(n9574), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[14] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14790.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14791 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[31] ), .I1(\lcd_data[15] ), 
            .I2(lcd_request), .O(n9575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14791.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14792 (.I0(n9575), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[15] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14792.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14793 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[32] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[16] ), 
            .I2(lcd_request), .O(n9576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14793.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14794 (.I0(n9576), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[16] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14794.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14795 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[33] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[17] ), 
            .I2(lcd_request), .O(n9577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14795.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14796 (.I0(n9577), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[17] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14796.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14797 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[34] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[18] ), 
            .I2(lcd_request), .O(n9578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14797.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14798 (.I0(n9578), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[18] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1489 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14798.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14799 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[35] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[19] ), 
            .I2(lcd_request), .O(n9579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14799.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14800 (.I0(n9579), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[19] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14800.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14801 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[36] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[20] ), 
            .I2(lcd_request), .O(n9580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14801.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14802 (.I0(n9580), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[20] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14802.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14803 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[37] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[21] ), 
            .I2(lcd_request), .O(n9581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14803.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14804 (.I0(n9581), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[21] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14804.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14805 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[38] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[22] ), 
            .I2(lcd_request), .O(n9582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14805.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14806 (.I0(n9582), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[22] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14806.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14807 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[39] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[23] ), 
            .I2(lcd_request), .O(n9583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14807.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14808 (.I0(n9583), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[23] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14808.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14809 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[40] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[24] ), 
            .I2(lcd_request), .O(n9584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14809.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14810 (.I0(n9584), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[24] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14810.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14811 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[41] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[25] ), 
            .I2(lcd_request), .O(n9585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14811.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14812 (.I0(n9585), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[25] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14812.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14813 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[42] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[26] ), 
            .I2(lcd_request), .O(n9586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14813.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14814 (.I0(n9586), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[26] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14814.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14815 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[43] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[27] ), 
            .I2(lcd_request), .O(n9587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14815.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14816 (.I0(n9587), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[27] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14816.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14817 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[44] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[28] ), 
            .I2(lcd_request), .O(n9588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14817.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14818 (.I0(n9588), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[28] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14818.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14819 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[45] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[29] ), 
            .I2(lcd_request), .O(n9589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14819.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14820 (.I0(n9589), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[29] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14820.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14821 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[46] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[30] ), 
            .I2(lcd_request), .O(n9590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14821.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14822 (.I0(n9590), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[30] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14822.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14823 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[47] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[31] ), 
            .I2(lcd_request), .O(n9591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14823.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14824 (.I0(n9591), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[31] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14824.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14825 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[48] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[32] ), 
            .I2(lcd_request), .O(n9592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14825.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14826 (.I0(n9592), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[32] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14826.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14827 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[49] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[33] ), 
            .I2(lcd_request), .O(n9593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14827.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14828 (.I0(n9593), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[33] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14828.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14829 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[50] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[34] ), 
            .I2(lcd_request), .O(n9594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14829.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14830 (.I0(n9594), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[34] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14830.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14831 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[51] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[35] ), 
            .I2(lcd_request), .O(n9595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14831.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14832 (.I0(n9595), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[35] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14832.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14833 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[52] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[36] ), 
            .I2(lcd_request), .O(n9596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14833.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14834 (.I0(n9596), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[36] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14834.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14835 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[53] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[37] ), 
            .I2(lcd_request), .O(n9597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14835.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14836 (.I0(n9597), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[37] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14836.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14837 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[54] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[38] ), 
            .I2(lcd_request), .O(n9598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14837.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14838 (.I0(n9598), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[38] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14838.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14839 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[55] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[39] ), 
            .I2(lcd_request), .O(n9599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14839.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14840 (.I0(n9599), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[39] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14840.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14841 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[56] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[40] ), 
            .I2(lcd_request), .O(n9600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14841.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14842 (.I0(n9600), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[40] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14842.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14843 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[57] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[41] ), 
            .I2(lcd_request), .O(n9601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14843.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14844 (.I0(n9601), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[41] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14844.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14845 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[58] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[42] ), 
            .I2(lcd_request), .O(n9602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14845.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14846 (.I0(n9602), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[42] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14846.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14847 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[59] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[43] ), 
            .I2(lcd_request), .O(n9603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14847.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14848 (.I0(n9603), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[43] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14848.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14849 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[60] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[44] ), 
            .I2(lcd_request), .O(n9604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14849.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14850 (.I0(n9604), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[44] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14850.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14851 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[61] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[45] ), 
            .I2(lcd_request), .O(n9605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14851.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14852 (.I0(n9605), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[45] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14852.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14853 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[62] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[46] ), 
            .I2(lcd_request), .O(n9606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14853.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14854 (.I0(n9606), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[46] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14854.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14855 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[63] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[47] ), 
            .I2(lcd_request), .O(n9607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14855.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14856 (.I0(n9607), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[47] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14856.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14857 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[64] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[48] ), 
            .I2(lcd_request), .O(n9608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14857.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14858 (.I0(n9608), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[48] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14858.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14859 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[65] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[49] ), 
            .I2(lcd_request), .O(n9609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14859.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14860 (.I0(n9609), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[49] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14860.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14861 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[66] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[50] ), 
            .I2(lcd_request), .O(n9610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14861.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14862 (.I0(n9610), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[50] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14862.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14863 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[67] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[51] ), 
            .I2(lcd_request), .O(n9611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14863.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14864 (.I0(n9611), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[51] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14864.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14865 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[68] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[52] ), 
            .I2(lcd_request), .O(n9612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14865.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14866 (.I0(n9612), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[52] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14866.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14867 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[69] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[53] ), 
            .I2(lcd_request), .O(n9613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14867.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14868 (.I0(n9613), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[53] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14868.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14869 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[70] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[54] ), 
            .I2(lcd_request), .O(n9614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14869.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14870 (.I0(n9614), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[54] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14870.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14871 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[71] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[55] ), 
            .I2(lcd_request), .O(n9615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14871.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14872 (.I0(n9615), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[55] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14872.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14873 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[72] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[56] ), 
            .I2(lcd_request), .O(n9616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14873.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14874 (.I0(n9616), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[56] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14874.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14875 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[73] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[57] ), 
            .I2(lcd_request), .O(n9617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14875.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14876 (.I0(n9617), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[57] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14876.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14877 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[74] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[58] ), 
            .I2(lcd_request), .O(n9618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14877.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14878 (.I0(n9618), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[58] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14878.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14879 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[75] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[59] ), 
            .I2(lcd_request), .O(n9619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14879.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14880 (.I0(n9619), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[59] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14880.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14881 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[76] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[60] ), 
            .I2(lcd_request), .O(n9620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14881.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14882 (.I0(n9620), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[60] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14882.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14883 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[77] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[61] ), 
            .I2(lcd_request), .O(n9621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14883.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14884 (.I0(n9621), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[61] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14884.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14885 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[78] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[62] ), 
            .I2(lcd_request), .O(n9622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14885.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14886 (.I0(n9622), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[62] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14886.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14887 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[79] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[63] ), 
            .I2(lcd_request), .O(n9623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14887.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14888 (.I0(n9623), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[63] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14888.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14889 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[80] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[64] ), 
            .I2(lcd_request), .O(n9624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14889.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14890 (.I0(n9624), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[64] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14890.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14891 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[81] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[65] ), 
            .I2(lcd_request), .O(n9625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14891.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14892 (.I0(n9625), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[65] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14892.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14893 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[82] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[66] ), 
            .I2(lcd_request), .O(n9626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14893.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14894 (.I0(n9626), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[66] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14894.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14895 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[83] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[67] ), 
            .I2(lcd_request), .O(n9627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14895.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14896 (.I0(n9627), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[67] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14896.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14897 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[84] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[68] ), 
            .I2(lcd_request), .O(n9628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14897.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14898 (.I0(n9628), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[68] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14898.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14899 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[85] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[69] ), 
            .I2(lcd_request), .O(n9629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14899.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14900 (.I0(n9629), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[69] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14900.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14901 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[86] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[70] ), 
            .I2(lcd_request), .O(n9630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14901.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14902 (.I0(n9630), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[70] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14902.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14903 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[87] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[71] ), 
            .I2(lcd_request), .O(n9631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14903.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14904 (.I0(n9631), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[71] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14904.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14905 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[88] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[72] ), 
            .I2(lcd_request), .O(n9632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14905.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14906 (.I0(n9632), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[72] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14906.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14907 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[89] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[73] ), 
            .I2(lcd_request), .O(n9633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14907.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14908 (.I0(n9633), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[73] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14908.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14909 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[90] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[74] ), 
            .I2(lcd_request), .O(n9634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14909.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14910 (.I0(n9634), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[74] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14910.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14911 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[91] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[75] ), 
            .I2(lcd_request), .O(n9635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14911.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14912 (.I0(n9635), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[75] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14912.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14913 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[92] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[76] ), 
            .I2(lcd_request), .O(n9636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14913.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14914 (.I0(n9636), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[76] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14914.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14915 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[93] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[77] ), 
            .I2(lcd_request), .O(n9637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14915.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14916 (.I0(n9637), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[77] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14916.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14917 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[94] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[78] ), 
            .I2(lcd_request), .O(n9638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14917.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14918 (.I0(n9638), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[78] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14918.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14919 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[95] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[79] ), 
            .I2(lcd_request), .O(n9639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14919.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14920 (.I0(n9639), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[79] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14920.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14921 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[96] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[80] ), 
            .I2(lcd_request), .O(n9640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14921.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14922 (.I0(n9640), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[80] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14922.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14923 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[97] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[81] ), 
            .I2(lcd_request), .O(n9641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14923.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14924 (.I0(n9641), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[81] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14924.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14925 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[98] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[82] ), 
            .I2(lcd_request), .O(n9642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14925.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14926 (.I0(n9642), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[82] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14926.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14927 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[99] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[83] ), 
            .I2(lcd_request), .O(n9643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14927.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14928 (.I0(n9643), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[83] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14928.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14929 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[100] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[84] ), 
            .I2(lcd_request), .O(n9644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14929.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14930 (.I0(n9644), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[84] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14930.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14931 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[101] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[85] ), 
            .I2(lcd_request), .O(n9645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14931.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14932 (.I0(n9645), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[85] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14932.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14933 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[102] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[86] ), 
            .I2(lcd_request), .O(n9646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14933.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14934 (.I0(n9646), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[86] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14934.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14935 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[103] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[87] ), 
            .I2(lcd_request), .O(n9647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14935.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14936 (.I0(n9647), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[87] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14936.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14937 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[104] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[88] ), 
            .I2(lcd_request), .O(n9648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14937.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14938 (.I0(n9648), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[88] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14938.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14939 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[105] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[89] ), 
            .I2(lcd_request), .O(n9649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14939.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14940 (.I0(n9649), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[89] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14940.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14941 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[106] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[90] ), 
            .I2(lcd_request), .O(n9650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14941.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14942 (.I0(n9650), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[90] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14942.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14943 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[107] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[91] ), 
            .I2(lcd_request), .O(n9651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14943.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14944 (.I0(n9651), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[91] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14944.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14945 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[108] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[92] ), 
            .I2(lcd_request), .O(n9652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14945.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14946 (.I0(n9652), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[92] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14946.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14947 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[109] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[93] ), 
            .I2(lcd_request), .O(n9653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14947.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14948 (.I0(n9653), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[93] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14948.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14949 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[110] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[94] ), 
            .I2(lcd_request), .O(n9654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14949.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14950 (.I0(n9654), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[94] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14950.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14951 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[111] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[95] ), 
            .I2(lcd_request), .O(n9655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14951.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14952 (.I0(n9655), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[95] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14952.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14953 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[112] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[96] ), 
            .I2(lcd_request), .O(n9656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14953.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14954 (.I0(n9656), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[96] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14954.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14955 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[113] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[97] ), 
            .I2(lcd_request), .O(n9657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14955.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14956 (.I0(n9657), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[97] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14956.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14957 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[114] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[98] ), 
            .I2(lcd_request), .O(n9658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14957.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14958 (.I0(n9658), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[98] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14958.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14959 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[115] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[99] ), 
            .I2(lcd_request), .O(n9659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14959.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14960 (.I0(n9659), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[99] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14960.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14961 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[116] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[100] ), 
            .I2(lcd_request), .O(n9660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14961.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14962 (.I0(n9660), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[100] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14962.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14963 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[117] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[101] ), 
            .I2(lcd_request), .O(n9661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14963.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14964 (.I0(n9661), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[101] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14964.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14965 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[118] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[102] ), 
            .I2(lcd_request), .O(n9662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14965.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14966 (.I0(n9662), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[102] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14966.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14967 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[119] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[103] ), 
            .I2(lcd_request), .O(n9663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14967.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14968 (.I0(n9663), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[103] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14968.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14969 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[120] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[104] ), 
            .I2(lcd_request), .O(n9664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14969.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14970 (.I0(n9664), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[104] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14970.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14971 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[121] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[105] ), 
            .I2(lcd_request), .O(n9665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14971.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14972 (.I0(n9665), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[105] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14972.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14973 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[122] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[106] ), 
            .I2(lcd_request), .O(n9666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14973.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14974 (.I0(n9666), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[106] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14974.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14975 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[123] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[107] ), 
            .I2(lcd_request), .O(n9667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14975.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14976 (.I0(n9667), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[107] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14976.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14977 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[124] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[108] ), 
            .I2(lcd_request), .O(n9668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14977.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14978 (.I0(n9668), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[108] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14978.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14979 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[125] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[109] ), 
            .I2(lcd_request), .O(n9669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14979.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14980 (.I0(n9669), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[109] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14980.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14981 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[126] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[110] ), 
            .I2(lcd_request), .O(n9670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14981.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14982 (.I0(n9670), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[110] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14982.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14983 (.I0(\u_axi4_ctrl_0/r_rframe_data_gen[127] ), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[111] ), 
            .I2(lcd_request), .O(n9671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__14983.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__14984 (.I0(n9671), .I1(\u_axi4_ctrl_0/w_rframe_data_gen[111] ), 
            .I2(n9544), .O(\u_axi4_ctrl_0/n1396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14984.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14985 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[112] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[112] ), .O(\u_axi4_ctrl_0/n1395 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14985.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14986 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[113] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[113] ), .O(\u_axi4_ctrl_0/n1394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14986.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14987 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[114] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[114] ), .O(\u_axi4_ctrl_0/n1393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14987.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14988 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[115] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[115] ), .O(\u_axi4_ctrl_0/n1392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14988.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14989 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[116] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[116] ), .O(\u_axi4_ctrl_0/n1391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14989.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14990 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[117] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[117] ), .O(\u_axi4_ctrl_0/n1390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14990.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14991 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[118] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[118] ), .O(\u_axi4_ctrl_0/n1389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14991.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14992 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[119] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[119] ), .O(\u_axi4_ctrl_0/n1388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14992.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14993 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[120] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[120] ), .O(\u_axi4_ctrl_0/n1387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14993.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14994 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[121] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[121] ), .O(\u_axi4_ctrl_0/n1386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14994.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14995 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[122] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[122] ), .O(\u_axi4_ctrl_0/n1385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14995.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14996 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[123] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[123] ), .O(\u_axi4_ctrl_0/n1384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14996.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14997 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[124] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[124] ), .O(\u_axi4_ctrl_0/n1383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14997.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14998 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[125] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[125] ), .O(\u_axi4_ctrl_0/n1382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14998.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__14999 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[126] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[126] ), .O(\u_axi4_ctrl_0/n1381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__14999.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15000 (.I0(lcd_request), .I1(\u_axi4_ctrl_0/r_rframe_data_gen[127] ), 
            .I2(n9544), .I3(\u_axi4_ctrl_0/w_rframe_data_gen[127] ), .O(\u_axi4_ctrl_0/n1380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15000.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15004 (.I0(DdrCtrl_ARREADY_0), .I1(DdrCtrl_ARVALID_0), 
            .I2(\DdrCtrl_ARADDR_0[8] ), .O(\u_axi4_ctrl_0/n1774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__15004.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__15005 (.I0(n1196), .I1(\DdrCtrl_ARADDR_0[9] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15005.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15006 (.I0(n631), .I1(\DdrCtrl_ARADDR_0[10] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15006.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15007 (.I0(n4368), .I1(\DdrCtrl_ARADDR_0[11] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15007.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15008 (.I0(n4366), .I1(\DdrCtrl_ARADDR_0[12] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15008.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15009 (.I0(n4364), .I1(\DdrCtrl_ARADDR_0[13] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15009.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15010 (.I0(n4362), .I1(\DdrCtrl_ARADDR_0[14] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15010.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15011 (.I0(n4360), .I1(\DdrCtrl_ARADDR_0[15] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15011.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15012 (.I0(n4358), .I1(\DdrCtrl_ARADDR_0[16] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15012.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15013 (.I0(n4356), .I1(\DdrCtrl_ARADDR_0[17] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15013.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15014 (.I0(n4354), .I1(\DdrCtrl_ARADDR_0[18] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15014.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15015 (.I0(n4352), .I1(\DdrCtrl_ARADDR_0[19] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15015.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15016 (.I0(n4350), .I1(\DdrCtrl_ARADDR_0[20] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15016.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15017 (.I0(n4349), .I1(\DdrCtrl_ARADDR_0[21] ), .I2(DdrCtrl_ARREADY_0), 
            .I3(DdrCtrl_ARVALID_0), .O(\u_axi4_ctrl_0/n1761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__15017.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__15021 (.I0(\DdrCtrl_ARADDR_0[22] ), .I1(n9531), .I2(\DdrCtrl_AWADDR_0[22] ), 
            .O(n9672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15021.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15022 (.I0(n9672), .I1(\u_axi4_ctrl_0/r_wframe_inc ), 
            .I2(\DdrCtrl_AWADDR_0[23] ), .O(\u_axi4_ctrl_0/n2772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__15022.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__15023 (.I0(\u_lcd_driver/vcnt[1] ), .I1(\u_lcd_driver/vcnt[0] ), 
            .I2(\u_lcd_driver/vcnt[2] ), .O(n9673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__15023.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__15024 (.I0(n9673), .I1(\u_lcd_driver/vcnt[3] ), .O(n9674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15024.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15025 (.I0(\u_lcd_driver/vcnt[5] ), .I1(\u_lcd_driver/vcnt[6] ), 
            .I2(\u_lcd_driver/vcnt[7] ), .O(n9675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15025.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15026 (.I0(n9674), .I1(\u_lcd_driver/vcnt[4] ), .I2(n9675), 
            .I3(\u_lcd_driver/vcnt[8] ), .O(n9676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__15026.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__15027 (.I0(\u_lcd_driver/vcnt[10] ), .I1(\u_lcd_driver/vcnt[11] ), 
            .O(n9677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15027.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15028 (.I0(\u_lcd_driver/hcnt[7] ), .I1(\u_lcd_driver/hcnt[8] ), 
            .I2(\u_lcd_driver/hcnt[11] ), .O(n9678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15028.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15029 (.I0(\u_lcd_driver/hcnt[2] ), .I1(\u_lcd_driver/hcnt[3] ), 
            .O(n9679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15029.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15030 (.I0(\u_lcd_driver/hcnt[0] ), .I1(\u_lcd_driver/hcnt[1] ), 
            .I2(n9679), .O(n9680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15030.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15031 (.I0(\u_lcd_driver/hcnt[4] ), .I1(\u_lcd_driver/hcnt[5] ), 
            .I2(\u_lcd_driver/hcnt[6] ), .O(n9681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15031.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15032 (.I0(\u_lcd_driver/hcnt[10] ), .I1(\u_lcd_driver/hcnt[9] ), 
            .I2(\u_lcd_driver/hcnt[11] ), .O(n9682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__15032.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__15033 (.I0(n9680), .I1(n9681), .I2(n9678), .I3(n9682), 
            .O(n9683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__15033.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__15034 (.I0(\u_lcd_driver/hcnt[1] ), .I1(n9678), .I2(n9679), 
            .I3(n9683), .O(n9684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15034.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15035 (.I0(\u_lcd_driver/vcnt[9] ), .I1(n9676), .I2(n9677), 
            .I3(n9684), .O(n9685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15035.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15036 (.I0(n9684), .I1(n9685), .I2(\u_lcd_driver/vcnt[0] ), 
            .O(\u_lcd_driver/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__15036.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__15037 (.I0(\u_lcd_driver/hcnt[3] ), .I1(\u_lcd_driver/hcnt[4] ), 
            .I2(\u_lcd_driver/hcnt[5] ), .I3(n9678), .O(n9686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__15037.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__15038 (.I0(\u_lcd_driver/hcnt[6] ), .I1(\u_lcd_driver/hcnt[9] ), 
            .I2(\u_lcd_driver/hcnt[10] ), .I3(n9686), .O(n9687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15038.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15039 (.I0(lcd_hs), .I1(n9687), .I2(r_hdmi_rst_n), .O(\u_lcd_driver/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__15039.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__15040 (.I0(\u_lcd_driver/vcnt[5] ), .I1(\u_lcd_driver/vcnt[6] ), 
            .I2(\u_lcd_driver/vcnt[7] ), .I3(\u_lcd_driver/vcnt[8] ), .O(n9688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15040.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15041 (.I0(\u_lcd_driver/vcnt[9] ), .I1(n9688), .O(n9689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15041.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15042 (.I0(n9673), .I1(\u_lcd_driver/vcnt[3] ), .I2(\u_lcd_driver/vcnt[4] ), 
            .I3(n9677), .O(n9690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15042.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15043 (.I0(n9690), .I1(n9689), .I2(lcd_vs), .I3(r_hdmi_rst_n), 
            .O(\u_lcd_driver/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__15043.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__15044 (.I0(\u_lcd_driver/hcnt[4] ), .I1(\u_lcd_driver/hcnt[5] ), 
            .I2(\u_lcd_driver/hcnt[6] ), .I3(\u_lcd_driver/hcnt[7] ), .O(n9691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15044.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15045 (.I0(n9679), .I1(n9691), .O(n9692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15045.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15046 (.I0(\u_lcd_driver/hcnt[9] ), .I1(n9692), .I2(\u_lcd_driver/hcnt[8] ), 
            .I3(\u_lcd_driver/hcnt[10] ), .O(n9693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5dba */ ;
    defparam LUT__15046.LUTMASK = 16'h5dba;
    EFX_LUT4 LUT__15047 (.I0(\u_lcd_driver/vcnt[0] ), .I1(\u_lcd_driver/vcnt[1] ), 
            .I2(\u_lcd_driver/vcnt[2] ), .I3(\u_lcd_driver/vcnt[3] ), .O(n9694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__15047.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__15048 (.I0(n9694), .I1(\u_lcd_driver/vcnt[4] ), .I2(n9675), 
            .I3(\u_lcd_driver/vcnt[8] ), .O(n9695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__15048.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__15049 (.I0(n9694), .I1(\u_lcd_driver/vcnt[4] ), .I2(n9689), 
            .I3(\u_lcd_driver/hcnt[11] ), .O(n9696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__15049.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__15050 (.I0(\u_lcd_driver/vcnt[9] ), .I1(n9695), .I2(n9677), 
            .I3(n9696), .O(n9697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15050.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15051 (.I0(n9693), .I1(n9697), .O(\u_lcd_driver/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15051.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15052 (.I0(\u_lcd_driver/hcnt[1] ), .I1(n9692), .I2(\u_lcd_driver/hcnt[8] ), 
            .I3(\u_lcd_driver/hcnt[10] ), .O(n9698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb4f */ ;
    defparam LUT__15052.LUTMASK = 16'hfb4f;
    EFX_LUT4 LUT__15053 (.I0(n9698), .I1(\u_lcd_driver/hcnt[9] ), .I2(\u_lcd_driver/hcnt[10] ), 
            .I3(n9697), .O(\u_lcd_driver/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d00 */ ;
    defparam LUT__15053.LUTMASK = 16'h7d00;
    EFX_LUT4 LUT__15054 (.I0(n9683), .I1(\u_lcd_driver/hcnt[0] ), .O(\u_lcd_driver/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15054.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15055 (.I0(n9684), .I1(\u_lcd_driver/vcnt[1] ), .I2(n9685), 
            .I3(n1653), .O(\u_lcd_driver/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15055.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15056 (.I0(n9684), .I1(\u_lcd_driver/vcnt[2] ), .I2(n9685), 
            .I3(n4192), .O(\u_lcd_driver/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15056.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15057 (.I0(n9684), .I1(\u_lcd_driver/vcnt[3] ), .I2(n9685), 
            .I3(n4190), .O(\u_lcd_driver/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15057.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15058 (.I0(n9684), .I1(\u_lcd_driver/vcnt[4] ), .I2(n9685), 
            .I3(n4188), .O(\u_lcd_driver/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15058.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15059 (.I0(n9684), .I1(\u_lcd_driver/vcnt[5] ), .I2(n9685), 
            .I3(n4186), .O(\u_lcd_driver/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15059.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15060 (.I0(n9684), .I1(\u_lcd_driver/vcnt[6] ), .I2(n9685), 
            .I3(n4184), .O(\u_lcd_driver/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15060.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15061 (.I0(n9684), .I1(\u_lcd_driver/vcnt[7] ), .I2(n9685), 
            .I3(n4182), .O(\u_lcd_driver/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15061.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15062 (.I0(n9684), .I1(\u_lcd_driver/vcnt[8] ), .I2(n9685), 
            .I3(n4180), .O(\u_lcd_driver/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15062.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15063 (.I0(n9684), .I1(\u_lcd_driver/vcnt[9] ), .I2(n9685), 
            .I3(n4178), .O(\u_lcd_driver/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15063.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15064 (.I0(n9684), .I1(\u_lcd_driver/vcnt[10] ), .I2(n9685), 
            .I3(n4176), .O(\u_lcd_driver/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15064.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15065 (.I0(n9684), .I1(\u_lcd_driver/vcnt[11] ), .I2(n9685), 
            .I3(n4175), .O(\u_lcd_driver/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__15065.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__15066 (.I0(n4556), .I1(n4558), .I2(n4560), .O(n9699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15066.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15067 (.I0(n4550), .I1(n4552), .I2(n4554), .O(n9700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15067.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15068 (.I0(n9699), .I1(n9700), .I2(n4548), .I3(n4547), 
            .O(n733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__15068.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__15069 (.I0(n9683), .I1(n1479), .O(\u_lcd_driver/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15069.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15070 (.I0(n9683), .I1(n4211), .O(\u_lcd_driver/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15070.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15071 (.I0(n9683), .I1(n4209), .O(\u_lcd_driver/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15071.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15072 (.I0(n9683), .I1(n4207), .O(\u_lcd_driver/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15072.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15073 (.I0(n9683), .I1(n4205), .O(\u_lcd_driver/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15073.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15074 (.I0(n9683), .I1(n4203), .O(\u_lcd_driver/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15074.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15075 (.I0(n9683), .I1(n4201), .O(\u_lcd_driver/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15075.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15076 (.I0(n9683), .I1(n4199), .O(\u_lcd_driver/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15076.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15077 (.I0(n9683), .I1(n4197), .O(\u_lcd_driver/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15077.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15078 (.I0(n9683), .I1(n4195), .O(\u_lcd_driver/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15078.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15079 (.I0(n9683), .I1(n4194), .O(\u_lcd_driver/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15079.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15080 (.I0(\u_lcd_driver/r_lcd_rgb[23] ), .I1(\u_lcd_driver/r_lcd_dv ), 
            .O(n9701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15080.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15081 (.I0(\u_black_pixel_avg/y_sum[0] ), .I1(n1716), 
            .I2(n9701), .O(\u_black_pixel_avg/n175 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15081.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15082 (.I0(n9701), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(\u_black_pixel_avg/n208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15082.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15083 (.I0(\u_black_pixel_avg/black_pixel_count[0] ), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .O(n9702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15083.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15084 (.I0(\u_black_pixel_avg/x_sum[27] ), .I1(n9702), 
            .O(n9703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15084.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15085 (.I0(\u_black_pixel_avg/x_sum[31] ), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .O(n9704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15085.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15086 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .O(n9705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15086.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15087 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[23] ), .I3(\u_black_pixel_avg/black_pixel_count[24] ), 
            .O(n9706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15087.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15088 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n9707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15088.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15089 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[12] ), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n9708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15089.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15090 (.I0(n9705), .I1(n9706), .I2(n9707), .I3(n9708), 
            .O(n9709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15090.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15091 (.I0(\u_black_pixel_avg/black_pixel_count[26] ), .I1(\u_black_pixel_avg/black_pixel_count[29] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[30] ), .I3(\u_black_pixel_avg/black_pixel_count[31] ), 
            .O(n9710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15091.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15092 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(\u_black_pixel_avg/black_pixel_count[25] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[27] ), .I3(\u_black_pixel_avg/black_pixel_count[28] ), 
            .O(n9711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15092.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15093 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n9712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15093.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15094 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .O(n9713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15094.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15095 (.I0(n9710), .I1(n9711), .I2(n9712), .I3(n9713), 
            .O(n9714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15095.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15096 (.I0(n9704), .I1(n9714), .I2(n9709), .I3(\u_black_pixel_avg/x_sum[30] ), 
            .O(n9715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__15096.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__15097 (.I0(\u_black_pixel_avg/x_sum[30] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15097.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15098 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n1812), 
            .I2(\u_black_pixel_avg/x_sum[31] ), .I3(n9716), .O(n9717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__15098.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__15099 (.I0(\u_black_pixel_avg/x_sum[30] ), .I1(n9702), 
            .I2(n1814), .O(n9718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15099.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15100 (.I0(n9717), .I1(n9714), .I2(n9709), .I3(n9718), 
            .O(n9719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15100.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15101 (.I0(n9715), .I1(n9719), .O(n6209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__15101.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__15102 (.I0(\u_black_pixel_avg/x_sum[29] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15102.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15103 (.I0(\u_black_pixel_avg/black_pixel_count[27] ), .I1(\u_black_pixel_avg/black_pixel_count[28] ), 
            .O(n9721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15103.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15104 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(\u_black_pixel_avg/black_pixel_count[25] ), 
            .O(n9722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15104.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15105 (.I0(n9721), .I1(n9710), .I2(n9722), .I3(n9706), 
            .O(n9723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15105.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15106 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .O(n9724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15106.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15107 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n9725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15107.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15108 (.I0(n9724), .I1(n9725), .I2(n9712), .O(n9726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15108.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15109 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n9727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15109.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15110 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[16] ), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n9728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15110.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15111 (.I0(n9727), .I1(n9728), .O(n9729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15111.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15112 (.I0(\u_black_pixel_avg/x_sum[31] ), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(\u_black_pixel_avg/x_sum[29] ), .I3(n9702), .O(n9730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15112.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15113 (.I0(n9723), .I1(n9726), .I2(n9729), .I3(n9730), 
            .O(n9731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15113.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15114 (.I0(n9720), .I1(n9719), .I2(n9715), .I3(n9731), 
            .O(n9732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__15114.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__15115 (.I0(\u_black_pixel_avg/x_sum[31] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15115.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15116 (.I0(n1812), .I1(n9714), .I2(n9733), .I3(n9709), 
            .O(n9734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15116.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15117 (.I0(n9709), .I1(n9714), .I2(n9733), .I3(\u_black_pixel_avg/x_sum[31] ), 
            .O(n9735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__15117.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__15118 (.I0(\u_black_pixel_avg/x_sum[30] ), .I1(n9702), 
            .I2(n1813), .O(n9736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15118.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15119 (.I0(n9736), .I1(n9714), .I2(n9709), .O(n9737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15119.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15120 (.I0(n9735), .I1(n9734), .I2(n9716), .I3(n9737), 
            .O(n9738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__15120.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__15121 (.I0(n6209), .I1(n1817), .I2(n9732), .I3(n9738), 
            .O(n6215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__15121.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__15122 (.I0(n6215), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n9739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15122.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15123 (.I0(\u_black_pixel_avg/x_sum[29] ), .I1(n1819), 
            .I2(n9732), .I3(n9738), .O(n6217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__15123.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__15124 (.I0(n6217), .I1(\u_black_pixel_avg/x_sum[28] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n9740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15124.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15125 (.I0(n9709), .I1(n9714), .O(n9741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15125.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15126 (.I0(n9736), .I1(\u_black_pixel_avg/x_sum[31] ), 
            .I2(n9709), .I3(n9714), .O(n9742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha333 */ ;
    defparam LUT__15126.LUTMASK = 16'ha333;
    EFX_LUT4 LUT__15127 (.I0(n9735), .I1(n9734), .I2(n9716), .I3(n9742), 
            .O(n6206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__15127.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__15128 (.I0(n9741), .I1(n1816), .I2(n9732), .I3(n6206), 
            .O(n6212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcdc0 */ ;
    defparam LUT__15128.LUTMASK = 16'hcdc0;
    EFX_LUT4 LUT__15129 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6215), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6212), .O(n9743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15129.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15130 (.I0(n9723), .I1(n9728), .O(n9744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15130.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15131 (.I0(n9744), .I1(n9726), .O(n9745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15131.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15132 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6212), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n9745), .O(n9746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15132.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15133 (.I0(n9739), .I1(n9740), .I2(n9743), .I3(n9746), 
            .O(n9747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15133.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15134 (.I0(\u_black_pixel_avg/x_sum[28] ), .I1(n1826), 
            .I2(n9703), .I3(n9747), .O(n9748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15134.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15135 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n1824), 
            .O(n9749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15135.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15136 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6217), 
            .O(n9750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15136.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15137 (.I0(\u_black_pixel_avg/x_sum[27] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15137.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15138 (.I0(n9750), .I1(n9749), .I2(n9751), .I3(n9747), 
            .O(n9752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__15138.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__15139 (.I0(n6215), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15139.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15140 (.I0(n6217), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n9754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15140.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15141 (.I0(n1822), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n1824), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n9755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15141.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15142 (.I0(n9754), .I1(n9753), .I2(n9755), .I3(n9747), 
            .O(n9756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__15142.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__15143 (.I0(n1822), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n1821), .O(n9757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15143.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15144 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6215), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n6212), .O(n9758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15144.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15145 (.I0(n9758), .I1(n9757), .I2(n9747), .O(n9759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15145.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15146 (.I0(n9748), .I1(n9752), .I2(n9756), .I3(n9759), 
            .O(n9760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15146.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15147 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6212), 
            .I2(n9745), .O(n9761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15147.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15148 (.I0(n1835), .I1(\u_black_pixel_avg/x_sum[27] ), 
            .I2(n9760), .I3(n9761), .O(n6239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15148.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15149 (.I0(n6217), .I1(n1824), .I2(n9747), .O(n6225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15149.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15150 (.I0(n1831), .I1(n6225), .I2(n9760), .I3(n9761), 
            .O(n6235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15150.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15151 (.I0(n6235), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15151.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15152 (.I0(\u_black_pixel_avg/x_sum[28] ), .I1(n1826), 
            .I2(n9747), .O(n6227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15152.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15153 (.I0(n1833), .I1(n6227), .I2(n9760), .I3(n9761), 
            .O(n6237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15153.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15154 (.I0(\u_black_pixel_avg/x_sum[26] ), .I1(n9702), 
            .I2(\u_black_pixel_avg/x_sum[27] ), .O(n9763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15154.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15155 (.I0(\u_black_pixel_avg/x_sum[26] ), .I1(n9702), 
            .I2(n1835), .I3(n9761), .O(n9764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__15155.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__15156 (.I0(\u_black_pixel_avg/x_sum[26] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n9765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15156.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15157 (.I0(n9765), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(n9761), .I3(\u_black_pixel_avg/x_sum[27] ), .O(n9766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8ee */ ;
    defparam LUT__15157.LUTMASK = 16'he8ee;
    EFX_LUT4 LUT__15158 (.I0(n9764), .I1(n9763), .I2(n9760), .I3(n9766), 
            .O(n9767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15158.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15159 (.I0(n6237), .I1(n9767), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n9768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4 */ ;
    defparam LUT__15159.LUTMASK = 16'hd4d4;
    EFX_LUT4 LUT__15160 (.I0(n6215), .I1(n1822), .I2(n9747), .O(n6223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15160.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15161 (.I0(n1829), .I1(n6223), .I2(n9760), .I3(n9761), 
            .O(n6233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15161.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15162 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6233), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6235), .O(n9769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15162.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15163 (.I0(n6212), .I1(n1821), .I2(n9747), .O(n6220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15163.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15164 (.I0(n1828), .I1(n6220), .I2(n9760), .I3(n9761), 
            .O(n6230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15164.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15165 (.I0(n6233), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n6230), .I3(\u_black_pixel_avg/black_pixel_count[5] ), .O(n9770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15165.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15166 (.I0(n9768), .I1(n9762), .I2(n9769), .I3(n9770), 
            .O(n9771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__15166.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__15167 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6230), 
            .O(n9772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15167.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15168 (.I0(n9709), .I1(n9710), .I2(n9711), .O(n9773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15168.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15169 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n9773), .O(n9774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15169.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15170 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n9774), 
            .O(n9775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15170.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15171 (.I0(n9772), .I1(n9771), .I2(n9775), .O(n9776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__15171.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__15172 (.I0(n6239), .I1(n1844), .I2(n9776), .O(n6251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15172.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15173 (.I0(n9772), .I1(n9771), .I2(n9775), .I3(n1846), 
            .O(n9777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__15173.LUTMASK = 16'he000;
    EFX_LUT4 LUT__15174 (.I0(\u_black_pixel_avg/x_sum[25] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15174.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15175 (.I0(n9772), .I1(n9771), .I2(n9775), .I3(\u_black_pixel_avg/x_sum[26] ), 
            .O(n9779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__15175.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__15176 (.I0(\u_black_pixel_avg/x_sum[25] ), .I1(n9702), 
            .O(n9780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15176.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15177 (.I0(n9778), .I1(n9779), .I2(n9777), .I3(n9780), 
            .O(n9781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__15177.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__15178 (.I0(n6237), .I1(n1842), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n9776), .O(n9782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15178.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15179 (.I0(n6251), .I1(n9781), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n9782), .O(n9783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__15179.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__15180 (.I0(n6237), .I1(n1842), .I2(n9776), .O(n6249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15180.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15181 (.I0(n6235), .I1(n1840), .I2(n9776), .O(n6247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15181.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15182 (.I0(n6247), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n6249), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n9784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15182.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15183 (.I0(n6233), .I1(n1838), .I2(n9776), .O(n6245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15183.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15184 (.I0(n6235), .I1(n1840), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n9776), .O(n9785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15184.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15185 (.I0(n6230), .I1(n1837), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n9776), .O(n9786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15185.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15186 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6245), 
            .I2(n9785), .I3(n9786), .O(n9787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__15186.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__15187 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6230), 
            .I2(n9774), .O(n9788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15187.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15188 (.I0(n6245), .I1(n9786), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n9788), .O(n9789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__15188.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__15189 (.I0(n9783), .I1(n9784), .I2(n9787), .I3(n9789), 
            .O(n9790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15189.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15190 (.I0(\u_black_pixel_avg/x_sum[25] ), .I1(n1859), 
            .I2(n9790), .O(n6269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15190.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15191 (.I0(n6230), .I1(n1837), .I2(n9776), .O(n6242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15191.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15192 (.I0(n6242), .I1(n1848), .I2(n9790), .O(n6256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15192.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15193 (.I0(\u_black_pixel_avg/x_sum[24] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(n1859), .O(n9791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15193.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15194 (.I0(\u_black_pixel_avg/x_sum[24] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/x_sum[25] ), 
            .O(n9792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15194.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15195 (.I0(\u_black_pixel_avg/x_sum[24] ), .I1(n9702), 
            .O(n9793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15195.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15196 (.I0(n9792), .I1(n9791), .I2(n9793), .I3(n9790), 
            .O(n9794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__15196.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__15197 (.I0(n9777), .I1(n9779), .O(n6253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__15197.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__15198 (.I0(n6253), .I1(n1857), .I2(n9790), .O(n6267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15198.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15199 (.I0(n6251), .I1(n1855), .I2(n9790), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15199.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15200 (.I0(n9794), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n6267), .I3(n9795), .O(n9796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15200.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15201 (.I0(n6251), .I1(n1855), .I2(n9790), .O(n6265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15201.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15202 (.I0(n6249), .I1(n1853), .I2(n9790), .O(n6263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15202.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15203 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6263), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6265), .O(n9797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15203.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15204 (.I0(n6247), .I1(n1851), .I2(n9790), .O(n6261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15204.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15205 (.I0(n6261), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6263), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n9798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15205.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15206 (.I0(n6245), .I1(n1849), .I2(n9790), .O(n6259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15206.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15207 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6259), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6261), .O(n9799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15207.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15208 (.I0(n9796), .I1(n9797), .I2(n9798), .I3(n9799), 
            .O(n9800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15208.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15209 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6259), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n9773), .O(n9801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15209.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15210 (.I0(n6256), .I1(n9800), .I2(n9774), .I3(n9801), 
            .O(n9802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4d5f */ ;
    defparam LUT__15210.LUTMASK = 16'h4d5f;
    EFX_LUT4 LUT__15211 (.I0(n1872), .I1(n6269), .I2(n9802), .O(n6285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15211.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15212 (.I0(n1868), .I1(n6265), .I2(n9802), .O(n6281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15212.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15213 (.I0(n1870), .I1(n6267), .I2(n9802), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15213.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15214 (.I0(n1866), .I1(n6263), .I2(n9802), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n9804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15214.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15215 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6281), 
            .I2(n9803), .I3(n9804), .O(n9805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15215.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15216 (.I0(\u_black_pixel_avg/x_sum[23] ), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[0] ), .O(n9806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15216.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15217 (.I0(\u_black_pixel_avg/x_sum[23] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15217.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15218 (.I0(n1874), .I1(\u_black_pixel_avg/x_sum[24] ), 
            .I2(n9807), .I3(n9802), .O(n9808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__15218.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__15219 (.I0(n6285), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n9806), .I3(n9808), .O(n9809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hddd4 */ ;
    defparam LUT__15219.LUTMASK = 16'hddd4;
    EFX_LUT4 LUT__15220 (.I0(n1870), .I1(n6267), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n9802), .O(n9810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15220.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15221 (.I0(n6281), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n9810), .I3(n9804), .O(n9811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15221.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15222 (.I0(n1866), .I1(n6263), .I2(n9802), .O(n6279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15222.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15223 (.I0(n1864), .I1(n6261), .I2(n9802), .O(n6277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15223.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15224 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6277), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6279), .O(n9812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15224.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15225 (.I0(n9809), .I1(n9805), .I2(n9811), .I3(n9812), 
            .O(n9813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__15225.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__15226 (.I0(n1862), .I1(n6259), .I2(n9802), .O(n6275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15226.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15227 (.I0(n1861), .I1(n6256), .I2(n9802), .O(n6272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15227.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15228 (.I0(n6272), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n6275), .I3(\u_black_pixel_avg/black_pixel_count[7] ), .O(n9814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15228.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15229 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6277), 
            .I2(n9814), .O(n9815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15229.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15230 (.I0(n6272), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6275), .O(n9816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15230.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15231 (.I0(n9813), .I1(n9815), .I2(n9816), .I3(n9773), 
            .O(n9817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15231.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15232 (.I0(n6285), .I1(n1887), .I2(n9817), .O(n6303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15232.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15233 (.I0(n1874), .I1(\u_black_pixel_avg/x_sum[24] ), 
            .I2(n9802), .O(n6287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15233.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15234 (.I0(n6287), .I1(n1889), .I2(n9817), .O(n6305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15234.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15235 (.I0(\u_black_pixel_avg/x_sum[22] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n9818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15235.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15236 (.I0(n9773), .I1(n1891), .O(n9819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15236.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15237 (.I0(n9813), .I1(n9815), .I2(n9816), .I3(n9819), 
            .O(n9820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15237.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15238 (.I0(n9773), .I1(n9816), .I2(\u_black_pixel_avg/x_sum[23] ), 
            .O(n9821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15238.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15239 (.I0(n9813), .I1(n9815), .I2(n9773), .I3(n9821), 
            .O(n9822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__15239.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__15240 (.I0(n9818), .I1(n9820), .I2(n9822), .I3(\u_black_pixel_avg/black_pixel_count[1] ), 
            .O(n9823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h54fd */ ;
    defparam LUT__15240.LUTMASK = 16'h54fd;
    EFX_LUT4 LUT__15241 (.I0(n6285), .I1(n1887), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n9817), .O(n9824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15241.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15242 (.I0(n6305), .I1(n9823), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n9824), .O(n9825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__15242.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__15243 (.I0(n1870), .I1(n6267), .I2(n9802), .O(n6283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15243.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15244 (.I0(n6283), .I1(n1885), .I2(n9817), .O(n6301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15244.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15245 (.I0(n6301), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n6303), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n9826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15245.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15246 (.I0(n6279), .I1(n1881), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n9817), .O(n9827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15246.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15247 (.I0(n6281), .I1(n1883), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n9817), .O(n9828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15247.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15248 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6301), 
            .I2(n9827), .I3(n9828), .O(n9829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__15248.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__15249 (.I0(n6279), .I1(n1881), .I2(n9817), .O(n6297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15249.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15250 (.I0(n6281), .I1(n1883), .I2(n9817), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n9830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15250.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15251 (.I0(n6277), .I1(n1879), .I2(n9817), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n9831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15251.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15252 (.I0(n6297), .I1(n9830), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n9831), .O(n9832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h002b */ ;
    defparam LUT__15252.LUTMASK = 16'h002b;
    EFX_LUT4 LUT__15253 (.I0(n9825), .I1(n9826), .I2(n9829), .I3(n9832), 
            .O(n9833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15253.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15254 (.I0(n6277), .I1(n1879), .I2(n9817), .O(n6295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15254.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15255 (.I0(n6275), .I1(n1877), .I2(n9817), .O(n6293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15255.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15256 (.I0(n6272), .I1(n1876), .I2(n9817), .O(n6290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15256.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15257 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6290), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6293), .O(n9834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15257.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15258 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6295), 
            .I2(n9834), .O(n9835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15258.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15259 (.I0(n6275), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .O(n9836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15259.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15260 (.I0(n9744), .I1(n9724), .O(n9837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15260.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15261 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n9837), 
            .O(n9838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15261.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15262 (.I0(n9836), .I1(n6290), .I2(n9838), .O(n9839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15262.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15263 (.I0(n6293), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n9773), .I3(n9839), .O(n9840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__15263.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__15264 (.I0(n9835), .I1(n9833), .I2(n9840), .O(n9841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15264.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15265 (.I0(n6303), .I1(n1904), .I2(n9841), .O(n6323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15265.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15266 (.I0(\u_black_pixel_avg/x_sum[22] ), .I1(n1910), 
            .I2(n9841), .O(n6329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15266.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15267 (.I0(\u_black_pixel_avg/x_sum[21] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n9842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15267.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15268 (.I0(n9822), .I1(n9820), .O(n6307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__15268.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__15269 (.I0(n6307), .I1(n1908), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n9841), .O(n9843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15269.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15270 (.I0(n6329), .I1(n9842), .I2(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I3(n9843), .O(n9844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__15270.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__15271 (.I0(n6301), .I1(n1902), .I2(n9841), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n9845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15271.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15272 (.I0(n6303), .I1(n1904), .I2(n9841), .I3(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n9846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15272.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15273 (.I0(n6305), .I1(n1906), .I2(n9841), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15273.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15274 (.I0(n6307), .I1(n1908), .I2(n9841), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n9848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15274.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15275 (.I0(n9845), .I1(n9846), .I2(n9847), .I3(n9848), 
            .O(n9849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15275.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15276 (.I0(n6305), .I1(n1906), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n9841), .O(n9850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15276.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15277 (.I0(n6323), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n9850), .I3(n9845), .O(n9851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15277.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15278 (.I0(n6301), .I1(n1902), .I2(n9841), .O(n6321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15278.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15279 (.I0(n6281), .I1(n1883), .I2(n9817), .O(n6299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15279.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15280 (.I0(n6299), .I1(n1900), .I2(n9841), .O(n6319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15280.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15281 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6319), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6321), .O(n9852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15281.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15282 (.I0(n9849), .I1(n9844), .I2(n9851), .I3(n9852), 
            .O(n9853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15282.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15283 (.I0(n6293), .I1(n1894), .I2(n9841), .O(n6313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15283.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15284 (.I0(n6295), .I1(n1896), .I2(n9841), .O(n6315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15284.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15285 (.I0(n6315), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n6313), .I3(\u_black_pixel_avg/black_pixel_count[9] ), .O(n9854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15285.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15286 (.I0(n6297), .I1(n1898), .I2(n9841), .O(n6317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15286.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15287 (.I0(n6317), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6319), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n9855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15287.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15288 (.I0(n9854), .I1(n9855), .O(n9856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15288.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15289 (.I0(n6315), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6317), .O(n9857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15289.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15290 (.I0(n6290), .I1(n1893), .I2(n9841), .O(n6310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15290.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15291 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6310), 
            .O(n9858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15291.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15292 (.I0(n9857), .I1(n6313), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(n9858), .O(n9859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15292.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15293 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6290), 
            .I2(n9837), .O(n9860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15293.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15294 (.I0(n9853), .I1(n9856), .I2(n9859), .I3(n9860), 
            .O(n9861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15294.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15295 (.I0(n6323), .I1(n1923), .I2(n9861), .O(n6345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15295.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15296 (.I0(n6305), .I1(n1906), .I2(n9841), .O(n6325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15296.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15297 (.I0(n6325), .I1(n1925), .I2(n9861), .O(n6347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15297.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15298 (.I0(n6307), .I1(n1908), .I2(n9841), .O(n6327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15298.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15299 (.I0(n6327), .I1(n1927), .I2(n9861), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15299.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15300 (.I0(n6323), .I1(n1923), .I2(n9861), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n9863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15300.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15301 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6347), 
            .I2(n9862), .I3(n9863), .O(n9864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15301.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15302 (.I0(n6329), .I1(n1929), .I2(n9861), .O(n6351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15302.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15303 (.I0(\u_black_pixel_avg/x_sum[20] ), .I1(n9702), 
            .O(n9865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15303.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15304 (.I0(\u_black_pixel_avg/x_sum[21] ), .I1(n1931), 
            .I2(n9865), .I3(n9861), .O(n9866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15304.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15305 (.I0(\u_black_pixel_avg/x_sum[20] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15305.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15306 (.I0(n6351), .I1(n9866), .I2(n9867), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n9868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe */ ;
    defparam LUT__15306.LUTMASK = 16'ha8fe;
    EFX_LUT4 LUT__15307 (.I0(n6327), .I1(n1927), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n9861), .O(n9869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15307.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15308 (.I0(n6347), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n9869), .I3(n9863), .O(n9870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15308.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15309 (.I0(n6321), .I1(n1921), .I2(n9861), .O(n6343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15309.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15310 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6343), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6345), .O(n9871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15310.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15311 (.I0(n9868), .I1(n9864), .I2(n9870), .I3(n9871), 
            .O(n9872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__15311.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__15312 (.I0(n6319), .I1(n1919), .I2(n9861), .O(n6341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15312.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15313 (.I0(n6341), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6343), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n9873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15313.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15314 (.I0(n6315), .I1(n1915), .I2(n9861), .O(n6337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15314.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15315 (.I0(n6313), .I1(n1913), .I2(n9861), .O(n6335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15315.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15316 (.I0(n6335), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n6337), .I3(\u_black_pixel_avg/black_pixel_count[9] ), .O(n9874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15316.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15317 (.I0(n6317), .I1(n1917), .I2(n9861), .O(n6339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15317.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15318 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n9744), .O(n9875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15318.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15319 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6310), 
            .I2(n9875), .O(n9876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15319.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15320 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6339), 
            .I2(n9876), .O(n9877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15320.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15321 (.I0(n9873), .I1(n9874), .I2(n9877), .O(n9878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15321.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15322 (.I0(n6339), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6341), .O(n9879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15322.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15323 (.I0(n6335), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6337), .O(n9880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15323.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15324 (.I0(n9879), .I1(n9874), .I2(n9880), .I3(n9876), 
            .O(n9881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15324.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15325 (.I0(n6310), .I1(n1912), .I2(n9861), .O(n6332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15325.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15326 (.I0(n6332), .I1(n9837), .O(n9882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15326.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15327 (.I0(n9878), .I1(n9872), .I2(n9881), .I3(n9882), 
            .O(n9883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15327.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15328 (.I0(n1944), .I1(n6345), .I2(n9883), .O(n6369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15328.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15329 (.I0(\u_black_pixel_avg/x_sum[21] ), .I1(n1931), 
            .I2(n9861), .O(n6353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15329.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15330 (.I0(n1952), .I1(n6353), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n9883), .O(n9884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15330.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15331 (.I0(\u_black_pixel_avg/x_sum[19] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/x_sum[20] ), 
            .O(n9885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15331.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15332 (.I0(\u_black_pixel_avg/x_sum[19] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(n1954), .O(n9886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15332.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15333 (.I0(\u_black_pixel_avg/x_sum[19] ), .I1(n9702), 
            .O(n9887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15333.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15334 (.I0(n9886), .I1(n9885), .I2(n9887), .I3(n9883), 
            .O(n9888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__15334.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__15335 (.I0(n1950), .I1(n6351), .I2(n9883), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15335.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15336 (.I0(n6327), .I1(n1927), .I2(n9861), .O(n6349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15336.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15337 (.I0(n6349), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n6353), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n9890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15337.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15338 (.I0(n1948), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n1952), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n9891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15338.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15339 (.I0(n9891), .I1(n9890), .I2(n9883), .O(n9892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15339.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15340 (.I0(n9888), .I1(n9884), .I2(n9889), .I3(n9892), 
            .O(n9893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__15340.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__15341 (.I0(n1948), .I1(n6349), .I2(n9883), .O(n6373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15341.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15342 (.I0(n1950), .I1(n6351), .I2(n9883), .O(n6375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15342.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15343 (.I0(n6373), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6375), .O(n9894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15343.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15344 (.I0(n1938), .I1(n6339), .I2(n9883), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n9895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15344.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15345 (.I0(n1940), .I1(n6341), .I2(n9883), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n9896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15345.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15346 (.I0(n6335), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n6337), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n9897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15346.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15347 (.I0(n1934), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n1936), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n9898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15347.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15348 (.I0(n9898), .I1(n9897), .I2(n9883), .O(n9899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15348.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15349 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6332), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n9744), 
            .O(n9900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15349.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15350 (.I0(n9895), .I1(n9896), .I2(n9899), .I3(n9900), 
            .O(n9901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15350.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15351 (.I0(n1946), .I1(n6347), .I2(n9883), .O(n6371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15351.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15352 (.I0(n1944), .I1(n6345), .I2(n9883), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n9902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15352.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15353 (.I0(n1942), .I1(n6343), .I2(n9883), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n9903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15353.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15354 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6371), 
            .I2(n9902), .I3(n9903), .O(n9904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15354.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15355 (.I0(n9894), .I1(n9893), .I2(n9901), .I3(n9904), 
            .O(n9905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15355.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15356 (.I0(n1938), .I1(n6339), .I2(n9883), .O(n6363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15356.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15357 (.I0(n1936), .I1(n6337), .I2(n9883), .O(n6361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15357.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15358 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6361), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6363), .O(n9906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15358.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15359 (.I0(n1933), .I1(n6332), .I2(n9883), .O(n6356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15359.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15360 (.I0(n1934), .I1(n6335), .I2(n9883), .O(n6359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15360.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15361 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6359), 
            .I2(\u_black_pixel_avg/black_pixel_count[12] ), .I3(n6356), 
            .O(n9907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15361.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15362 (.I0(n9899), .I1(n9906), .I2(n9907), .I3(n9900), 
            .O(n9908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__15362.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__15363 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6369), .I3(n6371), .O(n9909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15363.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15364 (.I0(n1940), .I1(n6341), .I2(n9883), .O(n6365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15364.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15365 (.I0(n1942), .I1(n6343), .I2(n9883), .O(n6367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15365.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15366 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6367), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6365), .O(n9910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15366.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15367 (.I0(n9903), .I1(n9909), .I2(n9910), .I3(n9901), 
            .O(n9911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__15367.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__15368 (.I0(n9905), .I1(n9908), .I2(n9911), .O(n9912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15368.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15369 (.I0(n1967), .I1(n6369), .I2(n9912), .O(n6395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15369.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15370 (.I0(n1954), .I1(\u_black_pixel_avg/x_sum[20] ), 
            .I2(n9883), .O(n6379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15370.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15371 (.I0(n1977), .I1(n6379), .I2(n9912), .O(n6405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15371.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15372 (.I0(\u_black_pixel_avg/x_sum[18] ), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[0] ), .O(n9913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15372.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15373 (.I0(n1979), .I1(\u_black_pixel_avg/x_sum[19] ), 
            .I2(n9913), .I3(n9912), .O(n9914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15373.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15374 (.I0(\u_black_pixel_avg/x_sum[18] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15374.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15375 (.I0(n6405), .I1(n9914), .I2(n9915), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n9916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe */ ;
    defparam LUT__15375.LUTMASK = 16'ha8fe;
    EFX_LUT4 LUT__15376 (.I0(n1973), .I1(n6375), .I2(n9912), .O(n6401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15376.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15377 (.I0(n1971), .I1(n6373), .I2(n9912), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n9917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15377.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15378 (.I0(n1952), .I1(n6353), .I2(n9883), .O(n6377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15378.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15379 (.I0(n1975), .I1(n6377), .I2(n9912), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15379.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15380 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6401), 
            .I2(n9917), .I3(n9918), .O(n9919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15380.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15381 (.I0(n1975), .I1(n6377), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n9912), .O(n9920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15381.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15382 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n9920), 
            .I2(n9917), .I3(n6401), .O(n9921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15382.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15383 (.I0(n6371), .I1(n1969), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n9912), .O(n9922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__15383.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__15384 (.I0(n6373), .I1(n1971), .I2(n9912), .O(n9923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__15384.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__15385 (.I0(n6377), .I1(n1975), .I2(n9912), .I3(n9727), 
            .O(n9924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__15385.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__15386 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n9924), 
            .I2(n9923), .I3(n9922), .O(n9925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15386.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15387 (.I0(n9919), .I1(n9916), .I2(n9921), .I3(n9925), 
            .O(n9926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__15387.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__15388 (.I0(n1959), .I1(n6361), .I2(n9912), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n9927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15388.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15389 (.I0(n1961), .I1(n6363), .I2(n9912), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n9928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15389.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15390 (.I0(n1963), .I1(n6365), .I2(n9912), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n9929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15390.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15391 (.I0(n1965), .I1(n6367), .I2(n9912), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n9930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15391.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15392 (.I0(n9927), .I1(n9928), .I2(n9929), .I3(n9930), 
            .O(n9931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15392.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15393 (.I0(n1969), .I1(n6371), .I2(n9912), .O(n6397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15393.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15394 (.I0(n6397), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n6395), .I3(\u_black_pixel_avg/black_pixel_count[7] ), .O(n9932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15394.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15395 (.I0(n9931), .I1(n9932), .O(n9933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15395.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15396 (.I0(n1965), .I1(n6367), .I2(n9912), .O(n6393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15396.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15397 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6395), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6393), .O(n9934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15397.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15398 (.I0(n1961), .I1(n6363), .I2(n9912), .O(n6389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15398.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15399 (.I0(n1963), .I1(n6365), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(n9912), .O(n9935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15399.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15400 (.I0(n6389), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n9935), .I3(n9927), .O(n9936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15400.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15401 (.I0(n1959), .I1(n6361), .I2(n9912), .O(n6387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15401.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15402 (.I0(n1957), .I1(n6359), .I2(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I3(n9912), .O(n9937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15402.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15403 (.I0(n1956), .I1(n6356), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n9912), .O(n9938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15403.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15404 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6387), 
            .I2(n9937), .I3(n9938), .O(n9939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__15404.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__15405 (.I0(n9934), .I1(n9931), .I2(n9936), .I3(n9939), 
            .O(n9940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__15405.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__15406 (.I0(n1956), .I1(n6356), .I2(n9912), .O(n6382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15406.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15407 (.I0(n1957), .I1(n6359), .I2(n9912), .O(n6385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15407.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15408 (.I0(n6382), .I1(n6385), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[12] ), .O(n9941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15408.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15409 (.I0(n9941), .I1(n9744), .O(n9942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15409.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15410 (.I0(n9926), .I1(n9933), .I2(n9940), .I3(n9942), 
            .O(n9943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15410.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15411 (.I0(n6395), .I1(n1992), .I2(n9943), .O(n6423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15411.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15412 (.I0(n6397), .I1(n1994), .I2(n9943), .O(n6425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15412.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15413 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6423), .I3(n6425), .O(n9944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15413.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15414 (.I0(n6393), .I1(n1990), .I2(n9943), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n9945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15414.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15415 (.I0(n1986), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n1988), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n9946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15415.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15416 (.I0(n1963), .I1(n6365), .I2(n9912), .O(n6391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15416.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15417 (.I0(n6391), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n6389), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n9947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15417.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15418 (.I0(n9947), .I1(n9946), .I2(n9943), .O(n9948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15418.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15419 (.I0(n6391), .I1(n1988), .I2(n9943), .O(n6419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15419.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15420 (.I0(n6393), .I1(n1990), .I2(n9943), .O(n6421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15420.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15421 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6421), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n6419), 
            .O(n9949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15421.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15422 (.I0(n9945), .I1(n9944), .I2(n9949), .I3(n9948), 
            .O(n9950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__15422.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__15423 (.I0(n1971), .I1(n6373), .I2(n9912), .O(n6399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15423.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15424 (.I0(n6399), .I1(n1996), .I2(n9943), .O(n6427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15424.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15425 (.I0(n2000), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n9951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15425.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15426 (.I0(n2006), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .O(n9952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15426.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15427 (.I0(n2006), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(\u_black_pixel_avg/x_sum[17] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n9953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15427.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15428 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n9952), 
            .I2(n9953), .I3(n2004), .O(n9954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe */ ;
    defparam LUT__15428.LUTMASK = 16'ha8fe;
    EFX_LUT4 LUT__15429 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2000), 
            .O(n9955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15429.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15430 (.I0(n9954), .I1(n2002), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n9955), .O(n9956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15430.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15431 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n9951), 
            .I2(n9956), .I3(n1998), .O(n9957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe */ ;
    defparam LUT__15431.LUTMASK = 16'ha8fe;
    EFX_LUT4 LUT__15432 (.I0(n1975), .I1(n6377), .I2(n9912), .O(n6403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15432.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15433 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6403), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6405), .O(n9958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15433.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15434 (.I0(n1979), .I1(\u_black_pixel_avg/x_sum[19] ), 
            .I2(n9912), .O(n6407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15434.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15435 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(\u_black_pixel_avg/x_sum[18] ), 
            .I2(\u_black_pixel_avg/x_sum[17] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n9959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15435.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15436 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6407), 
            .I2(n9959), .O(n9960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__15436.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__15437 (.I0(n6405), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n9960), .I3(n9958), .O(n9961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__15437.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__15438 (.I0(n6401), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6403), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n9962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15438.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15439 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6401), 
            .I2(n9961), .I3(n9962), .O(n9963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15439.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15440 (.I0(n9963), .I1(n9957), .I2(n9943), .O(n9964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15440.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15441 (.I0(n6427), .I1(n9964), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n9965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__15441.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__15442 (.I0(n6395), .I1(n1992), .I2(n9943), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n9966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15442.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15443 (.I0(n6397), .I1(n1994), .I2(n9943), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n9967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15443.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15444 (.I0(n9945), .I1(n9966), .I2(n9967), .I3(n9948), 
            .O(n9968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15444.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15445 (.I0(n6382), .I1(n1981), .I2(n9943), .O(n6410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15445.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15446 (.I0(n6385), .I1(n1982), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n9943), .O(n9969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15446.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15447 (.I0(n6410), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n9969), .O(n9970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__15447.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__15448 (.I0(n6387), .I1(n1984), .I2(n9943), .O(n6415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15448.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15449 (.I0(n6389), .I1(n1986), .I2(n9943), .O(n6417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15449.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15450 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6417), 
            .I2(\u_black_pixel_avg/black_pixel_count[12] ), .I3(n6415), 
            .O(n9971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15450.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15451 (.I0(n9968), .I1(n9965), .I2(n9970), .I3(n9971), 
            .O(n9972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__15451.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__15452 (.I0(n1982), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n1984), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n9973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15452.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15453 (.I0(n6385), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n6387), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n9974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15453.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15454 (.I0(n9974), .I1(n9973), .I2(n9969), .I3(n9943), 
            .O(n9975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__15454.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__15455 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n9723), 
            .O(n9976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15455.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15456 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n9976), 
            .O(n9977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15456.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15457 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n9977), 
            .O(n9978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15457.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15458 (.I0(n9975), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n6410), .I3(n9978), .O(n9979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__15458.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__15459 (.I0(n9972), .I1(n9950), .I2(n9979), .O(n9980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15459.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15460 (.I0(n6423), .I1(n2019), .I2(n9980), .O(n6453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15460.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15461 (.I0(\u_black_pixel_avg/x_sum[16] ), .I1(n9702), 
            .I2(n2035), .O(n9981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15461.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15462 (.I0(\u_black_pixel_avg/x_sum[16] ), .I1(n9702), 
            .I2(\u_black_pixel_avg/x_sum[17] ), .O(n9982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15462.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15463 (.I0(\u_black_pixel_avg/x_sum[16] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n9983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15463.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15464 (.I0(n9982), .I1(n9981), .I2(n9983), .I3(n9980), 
            .O(n9984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__15464.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__15465 (.I0(n6407), .I1(n2004), .I2(n9943), .O(n6435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15465.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15466 (.I0(n2031), .I1(n6435), .I2(n9980), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n9985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53 */ ;
    defparam LUT__15466.LUTMASK = 16'hac53;
    EFX_LUT4 LUT__15467 (.I0(\u_black_pixel_avg/x_sum[18] ), .I1(n2006), 
            .I2(n9943), .O(n6437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15467.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15468 (.I0(n6437), .I1(n2033), .I2(n9980), .O(n6467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15468.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15469 (.I0(n9984), .I1(n6467), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n9985), .O(n9986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__15469.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__15470 (.I0(n6405), .I1(n2002), .I2(n9943), .O(n6433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15470.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15471 (.I0(n6433), .I1(n2029), .I2(n9980), .O(n6463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15471.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15472 (.I0(n6435), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[2] ), .I3(n6437), .O(n9987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15472.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15473 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n2031), .I3(n2033), .O(n9988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15473.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15474 (.I0(n9988), .I1(n9987), .I2(n9980), .O(n9989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__15474.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__15475 (.I0(n6463), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n9989), .O(n9990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15475.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15476 (.I0(n6401), .I1(n1998), .I2(n9943), .O(n6429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15476.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15477 (.I0(n6429), .I1(n2025), .I2(n9980), .O(n6459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15477.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15478 (.I0(n6459), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n6463), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n9991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15478.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15479 (.I0(n6427), .I1(n2023), .I2(n9980), .O(n6457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15479.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15480 (.I0(n6403), .I1(n2000), .I2(n9943), .O(n6431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15480.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15481 (.I0(n6431), .I1(n2027), .I2(n9980), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n9992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15481.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15482 (.I0(n2019), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n2021), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n9993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15482.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15483 (.I0(n6423), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n6425), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n9994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15483.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15484 (.I0(n9994), .I1(n9993), .I2(n9980), .O(n9995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15484.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15485 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6457), 
            .I2(n9992), .I3(n9995), .O(n9996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15485.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15486 (.I0(n9990), .I1(n9986), .I2(n9991), .I3(n9996), 
            .O(n9997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15486.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15487 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6457), 
            .I2(n9995), .O(n9998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15487.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15488 (.I0(n6431), .I1(n2027), .I2(n9980), .O(n6461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15488.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15489 (.I0(n6459), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6461), .O(n9999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15489.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15490 (.I0(n6427), .I1(n2023), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n9980), .O(n10000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15490.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15491 (.I0(n6425), .I1(n2021), .I2(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I3(n9980), .O(n10001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15491.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15492 (.I0(n10001), .I1(n10000), .I2(n9995), .O(n10002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__15492.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__15493 (.I0(n6423), .I1(n2019), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(n9980), .O(n10003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15493.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15494 (.I0(n6421), .I1(n2017), .I2(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I3(n9980), .O(n10004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15494.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15495 (.I0(n6419), .I1(n2015), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(n9980), .O(n10005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15495.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15496 (.I0(n6417), .I1(n2013), .I2(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I3(n9980), .O(n10006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15496.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15497 (.I0(n10003), .I1(n10004), .I2(n10005), .I3(n10006), 
            .O(n10007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15497.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15498 (.I0(n9999), .I1(n9998), .I2(n10002), .I3(n10007), 
            .O(n10008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__15498.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__15499 (.I0(n6419), .I1(n2015), .I2(n9980), .O(n6449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15499.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15500 (.I0(n6421), .I1(n2017), .I2(n9980), .O(n6451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15500.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15501 (.I0(n6449), .I1(n6451), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[10] ), .O(n10009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15501.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15502 (.I0(n6417), .I1(n2013), .I2(n9980), .O(n6447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15502.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15503 (.I0(n6415), .I1(n2011), .I2(n9980), .O(n6445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15503.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15504 (.I0(n6445), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n6447), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n10010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15504.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15505 (.I0(n6385), .I1(n1982), .I2(n9943), .O(n6413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15505.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15506 (.I0(n6413), .I1(n2009), .I2(n9980), .O(n6443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15506.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15507 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n6410), 
            .I2(n9977), .O(n10011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15507.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15508 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n6443), 
            .I2(n10011), .O(n10012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15508.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15509 (.I0(n10006), .I1(n10009), .I2(n10010), .I3(n10012), 
            .O(n10013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__15509.LUTMASK = 16'he000;
    EFX_LUT4 LUT__15510 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n6445), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n6443), 
            .O(n10014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15510.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15511 (.I0(n6410), .I1(n2008), .I2(n9980), .O(n6440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15511.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15512 (.I0(n6440), .I1(n9978), .I2(n10014), .I3(n10012), 
            .O(n10015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__15512.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__15513 (.I0(n9997), .I1(n10008), .I2(n10013), .I3(n10015), 
            .O(n10016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15513.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15514 (.I0(n2048), .I1(n6453), .I2(n10016), .O(n6485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15514.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15515 (.I0(n6435), .I1(n2031), .I2(n9980), .O(n6465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15515.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15516 (.I0(n2060), .I1(n6465), .I2(n10016), .I3(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n10017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15516.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15517 (.I0(n6463), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n10018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15517.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15518 (.I0(\u_black_pixel_avg/x_sum[17] ), .I1(n2035), 
            .I2(n9980), .O(n6469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15518.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15519 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(\u_black_pixel_avg/x_sum[16] ), 
            .I2(\u_black_pixel_avg/x_sum[15] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15519.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15520 (.I0(n6469), .I1(n10019), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__15520.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__15521 (.I0(n10020), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n6467), .O(n10021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__15521.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__15522 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6465), 
            .I2(n10021), .O(n10022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15522.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15523 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2066), 
            .I2(\u_black_pixel_avg/x_sum[15] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15523.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15524 (.I0(n10023), .I1(n2064), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__15524.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__15525 (.I0(n10024), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n2062), .O(n10025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__15525.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__15526 (.I0(n2060), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n10025), .O(n10026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15526.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15527 (.I0(n2058), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n10026), .O(n10027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15527.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15528 (.I0(n10022), .I1(n10018), .I2(n10027), .I3(n10016), 
            .O(n10028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__15528.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__15529 (.I0(n2058), .I1(n6463), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n10016), .O(n10029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15529.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15530 (.I0(n2056), .I1(n6461), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n10016), .O(n10030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15530.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15531 (.I0(n10028), .I1(n10017), .I2(n10029), .I3(n10030), 
            .O(n10031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__15531.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__15532 (.I0(n2056), .I1(n6461), .I2(n10016), .O(n6493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15532.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15533 (.I0(n2054), .I1(n6459), .I2(n10016), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n10032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15533.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15534 (.I0(n6425), .I1(n2021), .I2(n9980), .O(n6455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15534.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15535 (.I0(n6455), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n6457), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15535.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15536 (.I0(n2050), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n2052), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15536.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15537 (.I0(n10034), .I1(n10033), .I2(n10016), .O(n10035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15537.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15538 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6493), 
            .I2(n10032), .I3(n10035), .O(n10036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15538.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15539 (.I0(n2050), .I1(n6455), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(n10016), .O(n10037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15539.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15540 (.I0(n2048), .I1(n6453), .I2(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I3(n10016), .O(n10038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15540.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15541 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6459), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6457), .O(n10039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15541.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15542 (.I0(n10039), .I1(n10033), .I2(n10016), .O(n10040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15542.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15543 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n2052), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n2054), .O(n10041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15543.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15544 (.I0(n10016), .I1(n10041), .I2(n10034), .O(n10042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15544.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15545 (.I0(n10037), .I1(n10038), .I2(n10040), .I3(n10042), 
            .O(n10043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15545.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15546 (.I0(n2046), .I1(n6451), .I2(n10016), .O(n6483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15546.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15547 (.I0(n6483), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n6485), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n10044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15547.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15548 (.I0(n10031), .I1(n10036), .I2(n10043), .I3(n10044), 
            .O(n10045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15548.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15549 (.I0(n2037), .I1(n6440), .I2(n10016), .O(n6472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15549.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15550 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n6472), 
            .O(n10046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15550.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15551 (.I0(n2042), .I1(n6447), .I2(n10016), .O(n6479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15551.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15552 (.I0(n2044), .I1(n6449), .I2(n10016), .O(n6481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15552.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15553 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6481), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n6479), 
            .O(n10047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15553.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15554 (.I0(n6445), .I1(n2040), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I3(n10016), .O(n10048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__15554.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__15555 (.I0(n6443), .I1(n2038), .I2(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I3(n10016), .O(n10049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__15555.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__15556 (.I0(n6483), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n10049), .I3(n10048), .O(n10050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15556.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15557 (.I0(n10046), .I1(n10047), .I2(n10050), .O(n10051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15557.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15558 (.I0(n2038), .I1(n6443), .I2(n10016), .O(n6475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15558.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15559 (.I0(n2040), .I1(n6445), .I2(n10016), .O(n6477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15559.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15560 (.I0(n6477), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n6475), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n10052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15560.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15561 (.I0(n6479), .I1(n6481), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[12] ), .O(n10053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15561.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15562 (.I0(n6475), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n6477), 
            .O(n10054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15562.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15563 (.I0(n10053), .I1(n10052), .I2(n10046), .I3(n10054), 
            .O(n10055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__15563.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__15564 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n6440), 
            .I2(n9976), .O(n10056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15564.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15565 (.I0(n10051), .I1(n10045), .I2(n10055), .I3(n10056), 
            .O(n10057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15565.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15566 (.I0(n6485), .I1(n2079), .I2(n10057), .O(n6514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15566.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15567 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2099), 
            .I2(\u_black_pixel_avg/x_sum[14] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15567.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15568 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(\u_black_pixel_avg/x_sum[15] ), 
            .I2(\u_black_pixel_avg/x_sum[14] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15568.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15569 (.I0(n10059), .I1(n10058), .I2(n10057), .O(n10060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15569.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15570 (.I0(n2066), .I1(\u_black_pixel_avg/x_sum[16] ), 
            .I2(n10016), .O(n6503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15570.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15571 (.I0(n6503), .I1(n2097), .I2(n10057), .O(n6532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15571.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15572 (.I0(n2064), .I1(n6469), .I2(n10016), .O(n6501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15572.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15573 (.I0(n6501), .I1(n2095), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15573.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15574 (.I0(n10060), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n6532), .I3(n10061), .O(n10062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15574.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15575 (.I0(n2058), .I1(n6463), .I2(n10016), .O(n6495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15575.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15576 (.I0(n6495), .I1(n2089), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n10057), .O(n10063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15576.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15577 (.I0(n2060), .I1(n6465), .I2(n10016), .O(n6497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15577.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15578 (.I0(n6497), .I1(n2091), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n10057), .O(n10064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15578.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15579 (.I0(n6501), .I1(n2095), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n10057), .O(n10065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15579.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15580 (.I0(n2062), .I1(n6467), .I2(n10016), .O(n6499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15580.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15581 (.I0(n6499), .I1(n2093), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n10057), .O(n10066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15581.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15582 (.I0(n10063), .I1(n10064), .I2(n10065), .I3(n10066), 
            .O(n10067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15582.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15583 (.I0(n6497), .I1(n2091), .I2(n10057), .O(n6526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15583.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15584 (.I0(n6499), .I1(n2093), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n10068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15584.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15585 (.I0(n6526), .I1(n10068), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n10063), .O(n10069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__15585.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__15586 (.I0(n6495), .I1(n2089), .I2(n10057), .O(n6524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15586.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15587 (.I0(n6493), .I1(n2087), .I2(n10057), .O(n6522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15587.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15588 (.I0(n6522), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6524), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15588.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15589 (.I0(n10067), .I1(n10062), .I2(n10069), .I3(n10070), 
            .O(n10071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15589.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15590 (.I0(n2054), .I1(n6459), .I2(n10016), .O(n6491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15590.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15591 (.I0(n6491), .I1(n2085), .I2(n10057), .O(n6520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15591.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15592 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6522), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6520), .O(n10072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15592.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15593 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n2077), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n2079), 
            .O(n10073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15593.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15594 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6483), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n6485), 
            .O(n10074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15594.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15595 (.I0(n10074), .I1(n10073), .I2(n10057), .O(n10075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15595.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15596 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n2081), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n2083), .O(n10076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15596.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15597 (.I0(n2050), .I1(n6455), .I2(n10016), .O(n6487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15597.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15598 (.I0(n2052), .I1(n6457), .I2(n10016), .O(n6489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15598.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15599 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6489), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n6487), 
            .O(n10077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15599.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15600 (.I0(n10077), .I1(n10076), .I2(n10057), .O(n10078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15600.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15601 (.I0(n10075), .I1(n10078), .I2(n10072), .O(n10079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15601.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15602 (.I0(n6491), .I1(n2085), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n10080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15602.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15603 (.I0(n6489), .I1(n2083), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n10081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15603.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15604 (.I0(n10081), .I1(n10080), .I2(n10075), .I3(n10078), 
            .O(n10082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__15604.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__15605 (.I0(n6487), .I1(n2081), .I2(n10057), .O(n6516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15605.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15606 (.I0(n6485), .I1(n2079), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n10083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15606.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15607 (.I0(n6516), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n10083), .I3(n10075), .O(n10084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15607.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15608 (.I0(n6481), .I1(n2075), .I2(n10057), .O(n6510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15608.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15609 (.I0(n6483), .I1(n2077), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n10085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15609.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15610 (.I0(n6479), .I1(n2073), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n10086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15610.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15611 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n6510), 
            .I2(n10085), .I3(n10086), .O(n10087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15611.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15612 (.I0(n6475), .I1(n2069), .I2(n10057), .O(n8372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15612.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15613 (.I0(n6477), .I1(n2071), .I2(n10057), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n10088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15613.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15614 (.I0(n9721), .I1(n9710), .O(n10089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15614.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15615 (.I0(\u_black_pixel_avg/black_pixel_count[25] ), .I1(n9706), 
            .I2(n10089), .O(n10090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15615.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15616 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I2(n10090), .O(n10091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15616.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15617 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n6472), 
            .I2(\u_black_pixel_avg/black_pixel_count[18] ), .I3(n10091), 
            .O(n10092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15617.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15618 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n8372), 
            .I2(n10088), .I3(n10092), .O(n10093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15618.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15619 (.I0(n10082), .I1(n10084), .I2(n10087), .I3(n10093), 
            .O(n10094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15619.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15620 (.I0(n6477), .I1(n2071), .I2(n10057), .O(n6506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15620.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15621 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n6506), 
            .O(n10095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15621.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15622 (.I0(n6479), .I1(n2073), .I2(n10057), .O(n6508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15622.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15623 (.I0(n6508), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n6510), 
            .O(n10096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15623.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15624 (.I0(n6472), .I1(n2068), .I2(n10057), .I3(n9976), 
            .O(n10097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__15624.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__15625 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n10092), 
            .I2(n8372), .I3(n10097), .O(n10098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__15625.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__15626 (.I0(n10095), .I1(n10096), .I2(n10093), .I3(n10098), 
            .O(n10099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15626.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15627 (.I0(n10071), .I1(n10079), .I2(n10094), .I3(n10099), 
            .O(n10100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15627.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15628 (.I0(n2109), .I1(n6514), .I2(n10100), .O(n6541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15628.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15629 (.I0(\u_black_pixel_avg/x_sum[15] ), .I1(n2099), 
            .I2(n10057), .O(n6534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15629.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15630 (.I0(n2129), .I1(n6534), .I2(n10100), .O(n6561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15630.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15631 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(\u_black_pixel_avg/x_sum[14] ), 
            .I2(\u_black_pixel_avg/x_sum[13] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15631.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15632 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2131), 
            .I2(\u_black_pixel_avg/x_sum[13] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15632.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15633 (.I0(n10102), .I1(n10101), .I2(n10100), .O(n10103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15633.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15634 (.I0(n2123), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2125), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15634.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15635 (.I0(n2127), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n2129), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n10105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15635.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15636 (.I0(n6534), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n6532), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n10106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15636.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15637 (.I0(n6501), .I1(n2095), .I2(n10057), .O(n6530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15637.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15638 (.I0(n6499), .I1(n2093), .I2(n10057), .O(n6528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15638.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15639 (.I0(n6528), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6530), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15639.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15640 (.I0(n10106), .I1(n10107), .O(n10108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15640.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15641 (.I0(n10105), .I1(n10104), .I2(n10108), .I3(n10100), 
            .O(n10109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__15641.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__15642 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6561), 
            .I2(n10103), .I3(n10109), .O(n10110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15642.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15643 (.I0(n2121), .I1(n6526), .I2(n10100), .O(n6553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15643.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15644 (.I0(n2123), .I1(n6528), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n10100), .O(n10111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15644.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15645 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2125), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n2127), .O(n10112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15645.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15646 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6530), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6532), .O(n10113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15646.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15647 (.I0(n10113), .I1(n10107), .O(n10114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15647.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15648 (.I0(n10112), .I1(n10104), .I2(n10114), .I3(n10100), 
            .O(n10115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__15648.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__15649 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6553), 
            .I2(n10111), .I3(n10115), .O(n10116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__15649.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__15650 (.I0(n2111), .I1(n6516), .I2(n10100), .O(n6543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15650.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15651 (.I0(n6489), .I1(n2083), .I2(n10057), .O(n6518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15651.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15652 (.I0(n2113), .I1(n6518), .I2(n10100), .O(n6545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15652.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15653 (.I0(n6545), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n6543), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n10117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15653.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15654 (.I0(n2115), .I1(n6520), .I2(n10100), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n10118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15654.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15655 (.I0(n2117), .I1(n6522), .I2(n10100), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n10119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15655.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15656 (.I0(n2119), .I1(n6524), .I2(n10100), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n10120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15656.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15657 (.I0(n2121), .I1(n6526), .I2(n10100), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n10121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15657.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15658 (.I0(n10118), .I1(n10119), .I2(n10120), .I3(n10121), 
            .O(n10122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15658.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15659 (.I0(n10116), .I1(n10110), .I2(n10117), .I3(n10122), 
            .O(n10123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15659.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15660 (.I0(n2117), .I1(n6522), .I2(n10100), .O(n6549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15660.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15661 (.I0(n2119), .I1(n6524), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n10100), .O(n10124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15661.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15662 (.I0(n6549), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n10124), .I3(n10118), .O(n10125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15662.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15663 (.I0(n2115), .I1(n6520), .I2(n10100), .O(n6547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15663.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15664 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6545), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6547), .O(n10126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15664.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15665 (.I0(n2105), .I1(n6510), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I3(n10100), .O(n10127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15665.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15666 (.I0(n6483), .I1(n2077), .I2(n10057), .O(n6512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15666.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15667 (.I0(n2107), .I1(n6512), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n10100), .O(n10128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15667.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15668 (.I0(n2111), .I1(n6516), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(n10100), .O(n10129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15668.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15669 (.I0(n2109), .I1(n6514), .I2(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I3(n10100), .O(n10130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15669.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15670 (.I0(n10127), .I1(n10128), .I2(n10129), .I3(n10130), 
            .O(n10131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15670.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15671 (.I0(n10125), .I1(n10126), .I2(n10117), .I3(n10131), 
            .O(n10132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15671.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15672 (.I0(n2107), .I1(n6512), .I2(n10100), .O(n6539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15672.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15673 (.I0(n2109), .I1(n6514), .I2(n10100), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n10133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15673.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15674 (.I0(n6539), .I1(n10133), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n10127), .O(n10134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__15674.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__15675 (.I0(n6472), .I1(n2068), .I2(n10057), .O(n8370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15675.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15676 (.I0(n3951), .I1(n8370), .I2(n10100), .O(n8362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15676.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15677 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n8362), 
            .I2(n10091), .O(n10135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15677.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15678 (.I0(n3952), .I1(n8372), .I2(n10100), .O(n8364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15678.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15679 (.I0(n2101), .I1(n6506), .I2(n10100), .O(n8366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15679.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15680 (.I0(n8366), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I2(n8364), .I3(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n10136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15680.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15681 (.I0(n2103), .I1(n6508), .I2(n10100), .O(n8368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15681.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15682 (.I0(n2105), .I1(n6510), .I2(n10100), .O(n6537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15682.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15683 (.I0(n6537), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n8368), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n10137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15683.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15684 (.I0(n10134), .I1(n10135), .I2(n10136), .I3(n10137), 
            .O(n10138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15684.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15685 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n8368), 
            .I2(\u_black_pixel_avg/black_pixel_count[16] ), .I3(n8366), 
            .O(n10139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15685.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15686 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n8362), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n8364), 
            .O(n10140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15686.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15687 (.I0(n10139), .I1(n10136), .I2(n10140), .I3(n10135), 
            .O(n10141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15687.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15688 (.I0(n10123), .I1(n10132), .I2(n10138), .I3(n10141), 
            .O(n10142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__15688.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__15689 (.I0(n2137), .I1(n6541), .I2(n10142), .O(n6566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15689.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15690 (.I0(n2131), .I1(\u_black_pixel_avg/x_sum[14] ), 
            .I2(n10100), .O(n6563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15690.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15691 (.I0(n2159), .I1(n6563), .I2(n10142), .O(n6588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15691.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15692 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6588), 
            .O(n10143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15692.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15693 (.I0(n2161), .I1(\u_black_pixel_avg/x_sum[13] ), 
            .I2(n10142), .O(n6590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15693.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15694 (.I0(n6590), .I1(\u_black_pixel_avg/x_sum[12] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15694.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15695 (.I0(n2127), .I1(n6532), .I2(n10100), .O(n6559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15695.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15696 (.I0(n2155), .I1(n6559), .I2(n10142), .O(n6584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15696.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15697 (.I0(n2125), .I1(n6530), .I2(n10100), .O(n6557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15697.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15698 (.I0(n2153), .I1(n6557), .I2(n10142), .O(n6582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15698.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15699 (.I0(n6582), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6584), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15699.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15700 (.I0(n2157), .I1(n6561), .I2(n10142), .O(n6586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15700.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15701 (.I0(n6586), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n6588), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n10146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15701.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15702 (.I0(n10144), .I1(n10143), .I2(n10145), .I3(n10146), 
            .O(n10147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__15702.LUTMASK = 16'he000;
    EFX_LUT4 LUT__15703 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6586), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n6584), .O(n10148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15703.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15704 (.I0(n2123), .I1(n6528), .I2(n10100), .O(n6555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15704.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15705 (.I0(n2151), .I1(n6555), .I2(n10142), .O(n6580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15705.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15706 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6580), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6582), .O(n10149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15706.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15707 (.I0(n10148), .I1(n10145), .I2(n10149), .O(n10150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15707.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15708 (.I0(n2149), .I1(n6553), .I2(n10142), .O(n6578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15708.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15709 (.I0(n6578), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6580), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15709.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15710 (.I0(n2141), .I1(n6545), .I2(n10142), .O(n6570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15710.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15711 (.I0(n2139), .I1(n6543), .I2(n10142), .O(n6568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15711.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15712 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6568), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n6570), 
            .O(n10152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15712.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15713 (.I0(n2119), .I1(n6524), .I2(n10100), .O(n6551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15713.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15714 (.I0(n2147), .I1(n6551), .I2(n10142), .O(n6576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15714.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15715 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6576), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6578), .O(n10153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15715.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15716 (.I0(n2145), .I1(n6549), .I2(n10142), .O(n6574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15716.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15717 (.I0(n2143), .I1(n6547), .I2(n10142), .O(n6572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15717.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15718 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6572), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6574), .O(n10154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15718.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15719 (.I0(n10152), .I1(n10153), .I2(n10154), .O(n10155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15719.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15720 (.I0(n10147), .I1(n10150), .I2(n10151), .I3(n10155), 
            .O(n10156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15720.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15721 (.I0(n3945), .I1(n8364), .I2(n10142), .O(n8352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15721.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15722 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n8362), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(n10090), 
            .O(n10157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15722.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15723 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n8352), 
            .I2(n10157), .O(n10158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15723.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15724 (.I0(n6574), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n6576), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15724.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15725 (.I0(n6572), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n6570), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n10160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15725.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15726 (.I0(n10159), .I1(n10154), .I2(n10160), .I3(n10152), 
            .O(n10161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15726.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15727 (.I0(n3949), .I1(n8368), .I2(n10142), .O(n8356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15727.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15728 (.I0(n2133), .I1(n6537), .I2(n10142), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n10162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15728.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15729 (.I0(n3947), .I1(n8366), .I2(n10142), .I3(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n10163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15729.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15730 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n8356), 
            .I2(n10162), .I3(n10163), .O(n10164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15730.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15731 (.I0(n2135), .I1(n6539), .I2(n10142), .O(n8360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15731.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15732 (.I0(n6566), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n8360), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n10165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15732.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15733 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6568), 
            .I2(n10164), .I3(n10165), .O(n10166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15733.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15734 (.I0(n10161), .I1(n10166), .O(n10167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15734.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15735 (.I0(n8360), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n6566), 
            .O(n10168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15735.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15736 (.I0(n2133), .I1(n6537), .I2(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I3(n10142), .O(n10169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15736.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15737 (.I0(n8356), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I2(n10169), .I3(n10163), .O(n10170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15737.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15738 (.I0(n3947), .I1(n8366), .I2(n10142), .O(n8354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15738.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15739 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n8352), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n8354), 
            .O(n10171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15739.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15740 (.I0(n10168), .I1(n10164), .I2(n10170), .I3(n10171), 
            .O(n10172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__15740.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__15741 (.I0(n3944), .I1(n8362), .I2(n10142), .O(n8350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15741.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15742 (.I0(n8350), .I1(n10091), .I2(n10172), .I3(n10158), 
            .O(n10173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__15742.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__15743 (.I0(n10156), .I1(n10167), .I2(n10158), .I3(n10173), 
            .O(n10174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__15743.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__15744 (.I0(n2163), .I1(n6566), .I2(n10174), .O(n8346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15744.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15745 (.I0(n2189), .I1(\u_black_pixel_avg/x_sum[12] ), 
            .I2(n10174), .O(n6615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15745.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15746 (.I0(\u_black_pixel_avg/x_sum[11] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15746.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15747 (.I0(n2187), .I1(n6590), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n10174), .O(n10176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15747.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15748 (.I0(n6615), .I1(n10175), .I2(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I3(n10176), .O(n10177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__15748.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__15749 (.I0(n2183), .I1(n6586), .I2(n10174), .I3(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n10178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15749.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15750 (.I0(n2181), .I1(n6584), .I2(n10174), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n10179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15750.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15751 (.I0(n2185), .I1(n6588), .I2(n10174), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15751.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15752 (.I0(n2187), .I1(n6590), .I2(n10174), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15752.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15753 (.I0(n10178), .I1(n10179), .I2(n10180), .I3(n10181), 
            .O(n10182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15753.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15754 (.I0(n2183), .I1(n6586), .I2(n10174), .O(n6609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15754.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15755 (.I0(n2185), .I1(n6588), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n10174), .O(n10183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15755.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15756 (.I0(n6609), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n10183), .I3(n10179), .O(n10184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15756.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15757 (.I0(n2181), .I1(n6584), .I2(n10174), .O(n6607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15757.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15758 (.I0(n2179), .I1(n6582), .I2(n10174), .O(n6605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15758.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15759 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6605), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6607), .O(n10185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15759.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15760 (.I0(n10182), .I1(n10177), .I2(n10184), .I3(n10185), 
            .O(n10186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15760.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15761 (.I0(n2171), .I1(n6574), .I2(n10174), .O(n6597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15761.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15762 (.I0(n2169), .I1(n6572), .I2(n10174), .O(n6595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15762.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15763 (.I0(n6595), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n6597), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n10187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15763.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15764 (.I0(n2175), .I1(n6578), .I2(n10174), .O(n6601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15764.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15765 (.I0(n2173), .I1(n6576), .I2(n10174), .O(n6599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15765.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15766 (.I0(n6599), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n6601), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15766.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15767 (.I0(n2177), .I1(n6580), .I2(n10174), .O(n6603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15767.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15768 (.I0(n6603), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6605), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15768.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15769 (.I0(n10187), .I1(n10188), .I2(n10189), .O(n10190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15769.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15770 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6603), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6601), .O(n10191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15770.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15771 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6599), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n6597), 
            .O(n10192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15771.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15772 (.I0(n10191), .I1(n10188), .I2(n10192), .I3(n10187), 
            .O(n10193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15772.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15773 (.I0(n2133), .I1(n6537), .I2(n10142), .O(n8358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15773.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15774 (.I0(n3940), .I1(n8358), .I2(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I3(n10174), .O(n10194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15774.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15775 (.I0(n3938), .I1(n8356), .I2(n10174), .O(n8340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15775.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15776 (.I0(n3936), .I1(n8354), .I2(n10174), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n10195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15776.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15777 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n10194), 
            .I2(n8340), .I3(n10195), .O(n10196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__15777.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__15778 (.I0(n3933), .I1(n8350), .I2(n10174), .O(n8334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15778.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15779 (.I0(n3936), .I1(n8354), .I2(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I3(n10174), .O(n10197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15779.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15780 (.I0(n3934), .I1(n8352), .I2(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I3(n10174), .O(n10198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15780.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15781 (.I0(\u_black_pixel_avg/black_pixel_count[20] ), .I1(n8334), 
            .I2(n10197), .I3(n10198), .O(n10199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__15781.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__15782 (.I0(n3942), .I1(n8360), .I2(n10174), .O(n8344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15782.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15783 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n8344), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n8346), 
            .O(n10200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15783.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15784 (.I0(n2167), .I1(n6570), .I2(n10174), .O(n6593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15784.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15785 (.I0(n2169), .I1(n6572), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(n10174), .O(n10201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15785.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15786 (.I0(n2165), .I1(n6568), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n10174), .O(n10202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15786.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15787 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6593), 
            .I2(n10201), .I3(n10202), .O(n10203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__15787.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__15788 (.I0(n10196), .I1(n10199), .I2(n10200), .I3(n10203), 
            .O(n10204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15788.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15789 (.I0(n10190), .I1(n10186), .I2(n10193), .I3(n10204), 
            .O(n10205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15789.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15790 (.I0(n2165), .I1(n6568), .I2(n10174), .O(n8348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15790.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15791 (.I0(n8348), .I1(n6593), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[12] ), .O(n10206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15791.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15792 (.I0(n8346), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n10206), .I3(n10200), .O(n10207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15792.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15793 (.I0(n3940), .I1(n8358), .I2(n10174), .O(n8342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15793.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15794 (.I0(n8340), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n8342), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n10208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15794.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15795 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n8344), 
            .I2(n10195), .I3(n10208), .O(n10209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15795.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15796 (.I0(n10196), .I1(n10199), .O(n10210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15796.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15797 (.I0(n3934), .I1(n8352), .I2(n10174), .O(n8336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15797.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15798 (.I0(n8334), .I1(n8336), .I2(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[19] ), .O(n10211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15798.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15799 (.I0(n10211), .I1(n10090), .O(n10212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15799.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15800 (.I0(n10207), .I1(n10209), .I2(n10210), .I3(n10212), 
            .O(n10213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15800.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15801 (.I0(n3929), .I1(n8346), .I2(n10205), .I3(n10213), 
            .O(n8326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15801.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15802 (.I0(n2215), .I1(\u_black_pixel_avg/x_sum[11] ), 
            .I2(n10205), .I3(n10213), .O(n6638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15802.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15803 (.I0(n6638), .I1(\u_black_pixel_avg/x_sum[10] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15803.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15804 (.I0(n10205), .I1(n10213), .O(n10215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15804.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15805 (.I0(n6615), .I1(n2213), .I2(n10215), .O(n6636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15805.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15806 (.I0(n2185), .I1(n6588), .I2(n10174), .O(n6611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15806.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15807 (.I0(n2209), .I1(n6611), .I2(n10205), .I3(n10213), 
            .O(n6632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15807.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15808 (.I0(n2187), .I1(n6590), .I2(n10174), .O(n6613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15808.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15809 (.I0(n2211), .I1(n6613), .I2(n10205), .I3(n10213), 
            .O(n6634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15809.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15810 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6634), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n6632), .O(n10216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15810.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15811 (.I0(n10214), .I1(n6636), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n10216), .O(n10217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__15811.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__15812 (.I0(n6609), .I1(n2207), .I2(n10215), .O(n6630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15812.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15813 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2209), 
            .I2(n2211), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n10218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15813.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15814 (.I0(n6611), .I1(n6613), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n10219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15814.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15815 (.I0(n10219), .I1(n10218), .I2(n10215), .O(n10220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15815.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15816 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6630), 
            .I2(n10220), .O(n10221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15816.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15817 (.I0(n6607), .I1(n2205), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n10215), .O(n10222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15817.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15818 (.I0(n6609), .I1(n2207), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n10215), .O(n10223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15818.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15819 (.I0(n2199), .I1(n6601), .I2(n10205), .I3(n10213), 
            .O(n6622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15819.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15820 (.I0(n2197), .I1(n6599), .I2(n10205), .I3(n10213), 
            .O(n6620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15820.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15821 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6620), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6622), .O(n10224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15821.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15822 (.I0(n2203), .I1(n6605), .I2(n10205), .I3(n10213), 
            .O(n6626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15822.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15823 (.I0(n2201), .I1(n6603), .I2(n10205), .I3(n10213), 
            .O(n6624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15823.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15824 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6624), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6626), .O(n10225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15824.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15825 (.I0(n10222), .I1(n10223), .I2(n10224), .I3(n10225), 
            .O(n10226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15825.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15826 (.I0(n10221), .I1(n10217), .I2(n10226), .O(n10227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15826.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15827 (.I0(n6607), .I1(n2205), .I2(n10215), .O(n6628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15827.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15828 (.I0(n6626), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n10228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15828.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15829 (.I0(n6628), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n10228), .I3(n10225), .O(n10229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__15829.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__15830 (.I0(n6624), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n6622), .I3(\u_black_pixel_avg/black_pixel_count[9] ), .O(n10230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15830.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15831 (.I0(n6620), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n10231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15831.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15832 (.I0(n2195), .I1(n6597), .I2(n10205), .I3(n10213), 
            .O(n6618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15832.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15833 (.I0(n6618), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n10232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15833.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15834 (.I0(n2193), .I1(n6595), .I2(n10205), .I3(n10213), 
            .O(n8332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15834.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15835 (.I0(n2191), .I1(n6593), .I2(n10205), .I3(n10213), 
            .O(n8330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15835.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15836 (.I0(n8330), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n8332), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n10233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15836.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15837 (.I0(n3931), .I1(n8348), .I2(n10205), .I3(n10213), 
            .O(n8328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15837.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15838 (.I0(n8326), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n8328), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n10234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15838.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15839 (.I0(n10231), .I1(n10232), .I2(n10233), .I3(n10234), 
            .O(n10235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15839.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15840 (.I0(n10229), .I1(n10230), .I2(n10224), .I3(n10235), 
            .O(n10236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15840.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15841 (.I0(n8332), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n6618), 
            .O(n10237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15841.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15842 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n8328), 
            .O(n10238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15842.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15843 (.I0(n10237), .I1(n8330), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n10238), .O(n10239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15843.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15844 (.I0(n8334), .I1(n3918), .I2(n10215), .I3(n10090), 
            .O(n10240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__15844.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__15845 (.I0(n3925), .I1(n8342), .I2(n10205), .I3(n10213), 
            .O(n8322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15845.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15846 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n8322), 
            .O(n10241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15846.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15847 (.I0(n3927), .I1(n8344), .I2(n10205), .I3(n10213), 
            .O(n8324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15847.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15848 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n8324), 
            .O(n10242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15848.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15849 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n8326), 
            .O(n10243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15849.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15850 (.I0(n10240), .I1(n10241), .I2(n10242), .I3(n10243), 
            .O(n10244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15850.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15851 (.I0(n8340), .I1(n3923), .I2(n10215), .O(n8320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15851.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15852 (.I0(n3919), .I1(n8336), .I2(n10205), .I3(n10213), 
            .O(n8316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15852.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15853 (.I0(n3936), .I1(n8354), .I2(n10174), .O(n8338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15853.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15854 (.I0(n3921), .I1(n8338), .I2(n10205), .I3(n10213), 
            .O(n8318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__15854.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__15855 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n8318), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(n8316), 
            .O(n10245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15855.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15856 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n8320), 
            .I2(n10245), .O(n10246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15856.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15857 (.I0(n10234), .I1(n10239), .I2(n10244), .I3(n10246), 
            .O(n10247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15857.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15858 (.I0(n8322), .I1(n8324), .I2(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[16] ), .O(n10248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15858.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15859 (.I0(n8320), .I1(n10248), .I2(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I3(n10245), .O(n10249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__15859.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__15860 (.I0(\u_black_pixel_avg/black_pixel_count[24] ), .I1(\u_black_pixel_avg/black_pixel_count[25] ), 
            .I2(n10089), .O(n10250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15860.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15861 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(n10250), 
            .O(n10251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15861.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15862 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n8334), 
            .I2(\u_black_pixel_avg/black_pixel_count[22] ), .I3(n10251), 
            .O(n10252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15862.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15863 (.I0(n8316), .I1(n8318), .I2(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[19] ), .O(n10253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15863.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15864 (.I0(n10249), .I1(n10253), .I2(n10252), .I3(n10240), 
            .O(n10254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__15864.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__15865 (.I0(n10227), .I1(n10236), .I2(n10247), .I3(n10254), 
            .O(n10255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__15865.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__15866 (.I0(n8326), .I1(n3910), .I2(n10255), .O(n8302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15866.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15867 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2239), 
            .I2(\u_black_pixel_avg/x_sum[9] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15867.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15868 (.I0(n2237), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n10256), .O(n10257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15868.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15869 (.I0(n2235), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n10257), .O(n10258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15869.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15870 (.I0(n6636), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n10258), .I3(n10255), .O(n10259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__15870.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__15871 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(\u_black_pixel_avg/x_sum[10] ), 
            .I2(\u_black_pixel_avg/x_sum[9] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15871.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15872 (.I0(n6638), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n10255), .I3(n10260), .O(n10261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15872.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15873 (.I0(n6638), .I1(n2237), .I2(n10255), .O(n6657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15873.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15874 (.I0(n6657), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n10261), .I3(n10259), .O(n10262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__15874.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__15875 (.I0(n6636), .I1(n2235), .I2(n10255), .O(n6655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15875.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15876 (.I0(n6634), .I1(n2233), .I2(n10255), .O(n6653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15876.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15877 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6653), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6655), .O(n10263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15877.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15878 (.I0(n6632), .I1(n2231), .I2(n10255), .O(n6651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15878.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15879 (.I0(n6651), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6653), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15879.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15880 (.I0(n6630), .I1(n2229), .I2(n10255), .O(n6649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15880.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15881 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6649), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6651), .O(n10265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15881.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15882 (.I0(n10262), .I1(n10263), .I2(n10264), .I3(n10265), 
            .O(n10266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15882.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15883 (.I0(n6622), .I1(n2221), .I2(n10255), .O(n6641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15883.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15884 (.I0(n6620), .I1(n2219), .I2(n10255), .O(n8312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15884.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15885 (.I0(n8312), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n6641), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n10267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15885.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15886 (.I0(n6626), .I1(n2225), .I2(n10255), .O(n6645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15886.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15887 (.I0(n6624), .I1(n2223), .I2(n10255), .O(n6643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15887.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15888 (.I0(n6643), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n6645), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15888.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15889 (.I0(n6628), .I1(n2227), .I2(n10255), .O(n6647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15889.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15890 (.I0(n6647), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6649), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15890.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15891 (.I0(n10267), .I1(n10268), .I2(n10269), .O(n10270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15891.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15892 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6647), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6645), .O(n10271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15892.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15893 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6643), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n6641), 
            .O(n10272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15893.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15894 (.I0(n10271), .I1(n10268), .I2(n10272), .I3(n10267), 
            .O(n10273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15894.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15895 (.I0(n8332), .I1(n3916), .I2(n10255), .O(n8308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15895.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15896 (.I0(n8330), .I1(n3914), .I2(n10255), .O(n8306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15896.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15897 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n8306), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n8308), 
            .O(n10274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15897.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15898 (.I0(n8328), .I1(n3912), .I2(n10255), .O(n8304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15898.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15899 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n8302), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n8304), 
            .O(n10275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15899.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15900 (.I0(n6618), .I1(n2217), .I2(n10255), .O(n8310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15900.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15901 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n8310), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n8312), 
            .O(n10276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15901.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15902 (.I0(n10274), .I1(n10275), .I2(n10276), .O(n10277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15902.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15903 (.I0(n10270), .I1(n10266), .I2(n10273), .I3(n10277), 
            .O(n10278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15903.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15904 (.I0(n8310), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n8308), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n10279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15904.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15905 (.I0(n8304), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n8306), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n10280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15905.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15906 (.I0(n10279), .I1(n10274), .I2(n10280), .I3(n10275), 
            .O(n10281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15906.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15907 (.I0(n8318), .I1(n3902), .I2(n10255), .O(n8294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15907.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15908 (.I0(n8316), .I1(n3900), .I2(n10255), .O(n8292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15908.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15909 (.I0(n8292), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I2(n8294), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n10282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15909.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15910 (.I0(n8320), .I1(n3904), .I2(n10255), .O(n8296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15910.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15911 (.I0(n8322), .I1(n3906), .I2(n10255), .O(n8298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15911.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15912 (.I0(n8298), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n8296), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n10283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15912.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15913 (.I0(n10282), .I1(n10283), .O(n10284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15913.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15914 (.I0(n8324), .I1(n3908), .I2(n10255), .O(n8300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15914.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15915 (.I0(n8300), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n8302), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n10285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15915.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15916 (.I0(n10281), .I1(n10284), .I2(n10285), .O(n10286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15916.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15917 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n8298), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n8300), 
            .O(n10287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15917.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15918 (.I0(n8334), .I1(n3918), .I2(n10215), .O(n8314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15918.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15919 (.I0(n8314), .I1(n3899), .I2(n10255), .O(n8290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15919.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15920 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n8290), 
            .O(n10288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15920.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15921 (.I0(n8294), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[19] ), .I3(n8296), 
            .O(n10289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15921.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15922 (.I0(n10289), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I2(n8292), .O(n10290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__15922.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__15923 (.I0(n10287), .I1(n10284), .I2(n10288), .I3(n10290), 
            .O(n10291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__15923.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__15924 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n8290), 
            .I2(n10251), .O(n10292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15924.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15925 (.I0(n10278), .I1(n10286), .I2(n10291), .I3(n10292), 
            .O(n10293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15925.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15926 (.I0(n8302), .I1(n3887), .I2(n10293), .O(n8274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15926.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15927 (.I0(n6651), .I1(n2251), .I2(n10293), .O(n6668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15927.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15928 (.I0(n6653), .I1(n2253), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n10293), .O(n10294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15928.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15929 (.I0(\u_black_pixel_avg/x_sum[10] ), .I1(n2239), 
            .I2(n10255), .O(n6659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15929.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15930 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(\u_black_pixel_avg/x_sum[9] ), 
            .I2(\u_black_pixel_avg/x_sum[8] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15930.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15931 (.I0(n6659), .I1(n10295), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__15931.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__15932 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6655), 
            .O(n10297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15932.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15933 (.I0(n10296), .I1(n6657), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n10297), .O(n10298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15933.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15934 (.I0(n6653), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6655), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15934.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15935 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2261), 
            .I2(\u_black_pixel_avg/x_sum[8] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15935.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15936 (.I0(n2257), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15936.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15937 (.I0(n10300), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n2259), .I3(n10301), .O(n10302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__15937.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__15938 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2255), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n2257), .O(n10303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15938.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15939 (.I0(n2253), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2255), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15939.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15940 (.I0(n10303), .I1(n10302), .I2(n10304), .O(n10305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15940.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15941 (.I0(n10298), .I1(n10299), .I2(n10305), .I3(n10293), 
            .O(n10306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__15941.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__15942 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6668), 
            .I2(n10294), .I3(n10306), .O(n10307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__15942.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__15943 (.I0(n6649), .I1(n2249), .I2(n10293), .O(n6666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15943.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15944 (.I0(n6666), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6668), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15944.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15945 (.I0(n6647), .I1(n2247), .I2(n10293), .O(n6664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15945.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15946 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6664), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6666), .O(n10309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15946.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15947 (.I0(n6645), .I1(n2245), .I2(n10293), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n10310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15947.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15948 (.I0(n6643), .I1(n2243), .I2(n10293), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n10311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15948.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15949 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6664), 
            .I2(n10310), .I3(n10311), .O(n10312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15949.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15950 (.I0(n10307), .I1(n10308), .I2(n10309), .I3(n10312), 
            .O(n10313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15950.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15951 (.I0(n8308), .I1(n3893), .I2(n10293), .O(n8280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15951.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15952 (.I0(n8310), .I1(n3895), .I2(n10293), .O(n8282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15952.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15953 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n8282), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n8280), 
            .O(n10314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15953.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15954 (.I0(n6643), .I1(n2243), .I2(n10293), .O(n8288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15954.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15955 (.I0(n6645), .I1(n2245), .I2(n10293), .O(n6662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15955.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15956 (.I0(n8288), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6662), .O(n10315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__15956.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__15957 (.I0(n8312), .I1(n3897), .I2(n10293), .O(n8284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15957.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15958 (.I0(n6641), .I1(n2241), .I2(n10293), .O(n8286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15958.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15959 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n8286), 
            .I2(\u_black_pixel_avg/black_pixel_count[12] ), .I3(n8284), 
            .O(n10316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15959.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15960 (.I0(n10314), .I1(n10315), .I2(n10316), .O(n10317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15960.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15961 (.I0(n8284), .I1(n8286), .I2(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[11] ), .O(n10318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15961.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15962 (.I0(n10318), .I1(n10314), .O(n10319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15962.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15963 (.I0(n8306), .I1(n3891), .I2(n10293), .O(n8278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15963.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15964 (.I0(n8278), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n10320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15964.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15965 (.I0(n8298), .I1(n3883), .I2(n10293), .O(n8270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15965.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15966 (.I0(n8300), .I1(n3885), .I2(n10293), .O(n8272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15966.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15967 (.I0(n8272), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n8270), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n10321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15967.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15968 (.I0(n8280), .I1(n8282), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[13] ), .O(n10322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15968.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15969 (.I0(n8304), .I1(n3889), .I2(n10293), .O(n8276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15969.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15970 (.I0(n8274), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n8276), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n10323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15970.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15971 (.I0(n10320), .I1(n10321), .I2(n10322), .I3(n10323), 
            .O(n10324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15971.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15972 (.I0(n10317), .I1(n10313), .I2(n10319), .I3(n10324), 
            .O(n10325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__15972.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__15973 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n8276), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n8278), 
            .O(n10326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15973.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15974 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n8274), 
            .I2(\u_black_pixel_avg/black_pixel_count[18] ), .I3(n8272), 
            .O(n10327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15974.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15975 (.I0(n10326), .I1(n10323), .I2(n10327), .I3(n10321), 
            .O(n10328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15975.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15976 (.I0(n8290), .I1(n3876), .I2(n10293), .O(n8262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15976.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15977 (.I0(n8292), .I1(n3877), .I2(n10293), .O(n8264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15977.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15978 (.I0(n8294), .I1(n3879), .I2(n10293), .O(n8266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15978.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15979 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n8266), 
            .I2(\u_black_pixel_avg/black_pixel_count[22] ), .I3(n8264), 
            .O(n10329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15979.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15980 (.I0(n10251), .I1(n8262), .I2(n10329), .O(n10330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__15980.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__15981 (.I0(n8296), .I1(n3881), .I2(n10293), .O(n8268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15981.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15982 (.I0(\u_black_pixel_avg/black_pixel_count[20] ), .I1(n8268), 
            .I2(\u_black_pixel_avg/black_pixel_count[19] ), .I3(n8270), 
            .O(n10331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15982.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15983 (.I0(n10328), .I1(n10330), .I2(n10331), .O(n10332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15983.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15984 (.I0(n8268), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I2(n8266), .I3(\u_black_pixel_avg/black_pixel_count[21] ), 
            .O(n10333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15984.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15985 (.I0(n8262), .I1(n8264), .I2(\u_black_pixel_avg/black_pixel_count[23] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[22] ), .O(n10334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__15985.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__15986 (.I0(n10333), .I1(n10330), .I2(n10334), .I3(n10250), 
            .O(n10335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__15986.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__15987 (.I0(n10332), .I1(n10325), .I2(n10335), .O(n10336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15987.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15988 (.I0(n8274), .I1(n3860), .I2(n10336), .O(n8242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15988.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15989 (.I0(\u_black_pixel_avg/x_sum[9] ), .I1(n2261), 
            .I2(n10293), .O(n6678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15989.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15990 (.I0(n6678), .I1(n2279), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15990.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15991 (.I0(\u_black_pixel_avg/x_sum[7] ), .I1(n9702), 
            .I2(\u_black_pixel_avg/x_sum[8] ), .O(n10338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15991.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15992 (.I0(\u_black_pixel_avg/x_sum[7] ), .I1(n9702), 
            .I2(n2281), .O(n10339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15992.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15993 (.I0(n10332), .I1(n10325), .I2(n10335), .I3(n10339), 
            .O(n10340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__15993.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__15994 (.I0(\u_black_pixel_avg/x_sum[7] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15994.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15995 (.I0(n10338), .I1(n10336), .I2(n10340), .I3(n10341), 
            .O(n10342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__15995.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__15996 (.I0(n6657), .I1(n2257), .I2(n10293), .O(n6674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15996.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15997 (.I0(n6674), .I1(n2275), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n10336), .O(n10343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15997.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15998 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n2277), 
            .I2(\u_black_pixel_avg/black_pixel_count[2] ), .I3(n2279), .O(n10344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__15998.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__15999 (.I0(n6659), .I1(n2259), .I2(n10293), .O(n6676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15999.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16000 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6676), 
            .I2(\u_black_pixel_avg/black_pixel_count[2] ), .I3(n6678), .O(n10345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16000.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16001 (.I0(n10345), .I1(n10344), .I2(n10336), .O(n10346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16001.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16002 (.I0(n10342), .I1(n10337), .I2(n10343), .I3(n10346), 
            .O(n10347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__16002.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__16003 (.I0(n6674), .I1(n2275), .I2(n10336), .O(n6689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16003.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16004 (.I0(n6676), .I1(n2277), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16004.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16005 (.I0(n6655), .I1(n2255), .I2(n10293), .O(n6672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16005.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16006 (.I0(n6672), .I1(n2273), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n10349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16006.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16007 (.I0(n6689), .I1(n10348), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n10349), .O(n10350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h002b */ ;
    defparam LUT__16007.LUTMASK = 16'h002b;
    EFX_LUT4 LUT__16008 (.I0(n6664), .I1(n2265), .I2(n10336), .O(n8260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16008.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16009 (.I0(n6662), .I1(n2263), .I2(n10336), .O(n8258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16009.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16010 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n8258), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n8260), .O(n10351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16010.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16011 (.I0(n6672), .I1(n2273), .I2(n10336), .O(n6687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16011.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16012 (.I0(n6653), .I1(n2253), .I2(n10293), .O(n6670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16012.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16013 (.I0(n6670), .I1(n2271), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n10336), .O(n10352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16013.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16014 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n2267), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n2269), .O(n10353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16014.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16015 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6666), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6668), .O(n10354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16015.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16016 (.I0(n10354), .I1(n10353), .I2(n10336), .O(n10355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__16016.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__16017 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6687), 
            .I2(n10352), .I3(n10355), .O(n10356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__16017.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__16018 (.I0(n10350), .I1(n10347), .I2(n10351), .I3(n10356), 
            .O(n10357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__16018.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__16019 (.I0(n2269), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n2271), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16019.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16020 (.I0(n6668), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6670), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16020.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16021 (.I0(n10359), .I1(n10358), .I2(n10336), .O(n10360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__16021.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__16022 (.I0(n6666), .I1(n2267), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n10361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16022.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16023 (.I0(n6664), .I1(n2265), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n10362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16023.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16024 (.I0(n10360), .I1(n10355), .I2(n10361), .I3(n10362), 
            .O(n10363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16024.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16025 (.I0(n8282), .I1(n3868), .I2(n10336), .O(n8250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16025.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16026 (.I0(n8280), .I1(n3866), .I2(n10336), .O(n8248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16026.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16027 (.I0(n8248), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n8250), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n10364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16027.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16028 (.I0(n8288), .I1(n3874), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n10365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16028.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16029 (.I0(n3870), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n3872), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n10366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16029.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16030 (.I0(n8286), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n8284), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n10367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16030.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16031 (.I0(n10367), .I1(n10366), .I2(n10336), .O(n10368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__16031.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__16032 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n8258), 
            .I2(n10365), .I3(n10368), .O(n10369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16032.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16033 (.I0(n10363), .I1(n10351), .I2(n10364), .I3(n10369), 
            .O(n10370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__16033.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__16034 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n3872), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n3874), 
            .O(n10371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16034.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16035 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n8286), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n8288), 
            .O(n10372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16035.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16036 (.I0(n10372), .I1(n10371), .I2(n10336), .O(n10373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__16036.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__16037 (.I0(n8282), .I1(n3868), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I3(n10336), .O(n10374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16037.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16038 (.I0(n8284), .I1(n3870), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n10336), .O(n10375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16038.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16039 (.I0(n10373), .I1(n10368), .I2(n10374), .I3(n10375), 
            .O(n10376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16039.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16040 (.I0(n8270), .I1(n3856), .I2(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I3(n10336), .O(n10377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16040.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16041 (.I0(n8272), .I1(n3858), .I2(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I3(n10336), .O(n10378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16041.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16042 (.I0(n8274), .I1(n3860), .I2(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I3(n10336), .O(n10379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16042.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16043 (.I0(n8276), .I1(n3862), .I2(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I3(n10336), .O(n10380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16043.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16044 (.I0(n10377), .I1(n10378), .I2(n10379), .I3(n10380), 
            .O(n10381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16044.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16045 (.I0(n8278), .I1(n3864), .I2(n10336), .O(n8246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16045.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16046 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n8248), 
            .I2(\u_black_pixel_avg/black_pixel_count[16] ), .I3(n8246), 
            .O(n10382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16046.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16047 (.I0(n10376), .I1(n10364), .I2(n10381), .I3(n10382), 
            .O(n10383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__16047.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__16048 (.I0(n8276), .I1(n3862), .I2(n10336), .O(n8244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16048.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16049 (.I0(n8246), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I2(n8244), .I3(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n10384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16049.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16050 (.I0(n8272), .I1(n3858), .I2(n10336), .O(n8240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16050.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16051 (.I0(n8274), .I1(n3860), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n10385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16051.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16052 (.I0(n8240), .I1(n10385), .I2(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I3(n10377), .O(n10386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__16052.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__16053 (.I0(n8266), .I1(n3852), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n10387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16053.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16054 (.I0(n8270), .I1(n3856), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n10388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16054.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16055 (.I0(n8268), .I1(n3854), .I2(n10336), .I3(\u_black_pixel_avg/black_pixel_count[21] ), 
            .O(n10389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16055.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16056 (.I0(n3850), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .O(n10390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16056.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16057 (.I0(n8264), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .O(n10391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16057.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16058 (.I0(\u_black_pixel_avg/black_pixel_count[24] ), .I1(n8262), 
            .I2(\u_black_pixel_avg/black_pixel_count[25] ), .I3(n10089), 
            .O(n10392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__16058.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__16059 (.I0(n10391), .I1(n10390), .I2(n10336), .I3(n10392), 
            .O(n10393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16059.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16060 (.I0(n10387), .I1(n10388), .I2(n10389), .I3(n10393), 
            .O(n10394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__16060.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__16061 (.I0(n10384), .I1(n10381), .I2(n10386), .I3(n10394), 
            .O(n10395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__16061.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__16062 (.I0(n10357), .I1(n10370), .I2(n10383), .I3(n10395), 
            .O(n10396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16062.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16063 (.I0(n8262), .I1(n3849), .I2(n10336), .O(n8230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16063.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16064 (.I0(n8264), .I1(n3850), .I2(n10336), .O(n8232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16064.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16065 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(n8232), 
            .I2(\u_black_pixel_avg/black_pixel_count[24] ), .I3(n8230), 
            .O(n10397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16065.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16066 (.I0(n8266), .I1(n3852), .I2(n10336), .O(n8234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16066.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16067 (.I0(n8268), .I1(n3854), .I2(n10336), .O(n8236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16067.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16068 (.I0(n8234), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(n8236), 
            .O(n10398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16068.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16069 (.I0(n10398), .I1(n10393), .I2(n10397), .I3(n10392), 
            .O(n10399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16069.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16070 (.I0(n10396), .I1(n10399), .O(n10400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16070.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16071 (.I0(n3829), .I1(n8242), .I2(n10400), .O(n8206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16071.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16072 (.I0(n6678), .I1(n2279), .I2(n10336), .O(n6693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16072.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16073 (.I0(n6693), .I1(n2295), .I2(n10396), .I3(n10399), 
            .O(n6706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16073.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16074 (.I0(n6706), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16074.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16075 (.I0(\u_black_pixel_avg/x_sum[6] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16075.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16076 (.I0(n10402), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(\u_black_pixel_avg/x_sum[7] ), .O(n10403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__16076.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__16077 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n10403), 
            .O(n10404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16077.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16078 (.I0(n10402), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(n2299), .O(n10405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__16078.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__16079 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n10405), 
            .O(n10406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16079.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16080 (.I0(\u_black_pixel_avg/x_sum[8] ), .I1(n2281), 
            .I2(n10336), .O(n6695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16080.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16081 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n10403), 
            .I2(n6695), .O(n10407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16081.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16082 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n10405), 
            .I2(n2297), .O(n10408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16082.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16083 (.I0(n10407), .I1(n10408), .I2(n10396), .I3(n10399), 
            .O(n10409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__16083.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__16084 (.I0(n10406), .I1(n10404), .I2(n10400), .I3(n10409), 
            .O(n10410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16084.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16085 (.I0(n6676), .I1(n2277), .I2(n10336), .O(n6691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16085.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16086 (.I0(n6691), .I1(n2293), .I2(n10396), .I3(n10399), 
            .O(n6704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16086.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16087 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6704), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6706), .O(n10411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16087.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16088 (.I0(n6689), .I1(n2291), .I2(n10396), .I3(n10399), 
            .O(n6702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16088.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16089 (.I0(n6702), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6704), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16089.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16090 (.I0(n10410), .I1(n10401), .I2(n10411), .I3(n10412), 
            .O(n10413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__16090.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__16091 (.I0(n6687), .I1(n2289), .I2(n10396), .I3(n10399), 
            .O(n6700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16091.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16092 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6700), 
            .O(n10414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16092.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16093 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6702), 
            .O(n10415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16093.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16094 (.I0(n6666), .I1(n2267), .I2(n10336), .O(n6681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16094.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16095 (.I0(n6681), .I1(n2283), .I2(n10396), .I3(n10399), 
            .O(n8226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16095.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16096 (.I0(n8260), .I1(n3847), .I2(n10396), .I3(n10399), 
            .O(n8224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16096.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16097 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n8224), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n8226), .O(n10416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16097.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16098 (.I0(n6670), .I1(n2271), .I2(n10336), .O(n6685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16098.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16099 (.I0(n6685), .I1(n2287), .I2(n10396), .I3(n10399), 
            .O(n6698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16099.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16100 (.I0(n6668), .I1(n2269), .I2(n10336), .O(n6683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16100.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16101 (.I0(n6683), .I1(n2285), .I2(n10396), .I3(n10399), 
            .O(n8228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16101.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16102 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n8228), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6698), .O(n10417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16102.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16103 (.I0(n10414), .I1(n10415), .I2(n10416), .I3(n10417), 
            .O(n10418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__16103.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__16104 (.I0(n6700), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n6698), .I3(\u_black_pixel_avg/black_pixel_count[7] ), .O(n10419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16104.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16105 (.I0(n8228), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n8226), .I3(\u_black_pixel_avg/black_pixel_count[9] ), .O(n10420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16105.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16106 (.I0(n10419), .I1(n10417), .I2(n10420), .I3(n10416), 
            .O(n10421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16106.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16107 (.I0(n8224), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n10422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16107.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16108 (.I0(n3845), .I1(n8258), .I2(n10400), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n10423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16108.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16109 (.I0(n8250), .I1(n3837), .I2(n10396), .I3(n10399), 
            .O(n8214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16109.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16110 (.I0(n8284), .I1(n3870), .I2(n10336), .O(n8252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16110.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16111 (.I0(n8252), .I1(n3839), .I2(n10396), .I3(n10399), 
            .O(n8216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16111.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16112 (.I0(n8216), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n8214), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n10424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16112.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16113 (.I0(n8288), .I1(n3874), .I2(n10336), .O(n8256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16113.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16114 (.I0(n8256), .I1(n3843), .I2(n10396), .I3(n10399), 
            .O(n8220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16114.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16115 (.I0(n8286), .I1(n3872), .I2(n10336), .O(n8254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16115.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16116 (.I0(n8254), .I1(n3841), .I2(n10399), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n10425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__16116.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__16117 (.I0(n3841), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n10425), .I3(n10396), .O(n10426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__16117.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__16118 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n8220), 
            .I2(n10426), .O(n10427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16118.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16119 (.I0(n10422), .I1(n10423), .I2(n10424), .I3(n10427), 
            .O(n10428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__16119.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__16120 (.I0(n10418), .I1(n10413), .I2(n10421), .I3(n10428), 
            .O(n10429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__16120.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__16121 (.I0(n8254), .I1(n3841), .I2(n10396), .I3(n10399), 
            .O(n8218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16121.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16122 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n8218), 
            .O(n10430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16122.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16123 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n8216), 
            .O(n10431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16123.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16124 (.I0(n8258), .I1(n3845), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(n10399), .O(n10432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__16124.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__16125 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n3845), 
            .I2(n10432), .I3(n10396), .O(n10433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__16125.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__16126 (.I0(n8220), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n10433), .I3(n10426), .O(n10434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b00 */ ;
    defparam LUT__16126.LUTMASK = 16'h2b00;
    EFX_LUT4 LUT__16127 (.I0(n10431), .I1(n10434), .I2(n10430), .I3(n10424), 
            .O(n10435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__16127.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__16128 (.I0(n8232), .I1(n3819), .I2(n10396), .I3(n10399), 
            .O(n8196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16128.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16129 (.I0(n8234), .I1(n3821), .I2(n10396), .I3(n10399), 
            .O(n8198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16129.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16130 (.I0(n8198), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .I2(n8196), .I3(\u_black_pixel_avg/black_pixel_count[24] ), 
            .O(n10436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16130.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16131 (.I0(n8236), .I1(n3823), .I2(n10396), .I3(n10399), 
            .O(n8200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16131.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16132 (.I0(n8270), .I1(n3856), .I2(n10336), .O(n8238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16132.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16133 (.I0(n8238), .I1(n3825), .I2(n10396), .I3(n10399), 
            .O(n8202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16133.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16134 (.I0(n8200), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(n8202), 
            .O(n10437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16134.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16135 (.I0(n3818), .I1(n8230), .I2(\u_black_pixel_avg/black_pixel_count[25] ), 
            .I3(n10400), .O(n10438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16135.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16136 (.I0(n8196), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[23] ), .I3(n8198), 
            .O(n10439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16136.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16137 (.I0(n10437), .I1(n10436), .I2(n10438), .I3(n10439), 
            .O(n10440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__16137.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__16138 (.I0(n3827), .I1(n8240), .I2(n10400), .O(n8204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16138.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16139 (.I0(\u_black_pixel_avg/black_pixel_count[20] ), .I1(n8204), 
            .I2(\u_black_pixel_avg/black_pixel_count[19] ), .I3(n8206), 
            .O(n10441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16139.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16140 (.I0(n8248), .I1(n3835), .I2(n10396), .I3(n10399), 
            .O(n8212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16140.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16141 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n8214), 
            .O(n10442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16141.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16142 (.I0(n8246), .I1(n3833), .I2(n10396), .I3(n10399), 
            .O(n8210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16142.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16143 (.I0(n8244), .I1(n3831), .I2(n10396), .I3(n10399), 
            .O(n8208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__16143.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__16144 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n8208), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n8210), 
            .O(n10443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16144.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16145 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n8212), 
            .I2(n10442), .I3(n10443), .O(n10444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__16145.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__16146 (.I0(n10435), .I1(n10440), .I2(n10441), .I3(n10444), 
            .O(n10445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__16146.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__16147 (.I0(n8210), .I1(n8212), .I2(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[16] ), .O(n10446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16147.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16148 (.I0(n3829), .I1(n8242), .I2(n10400), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n10447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16148.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16149 (.I0(n10446), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n8208), .I3(n10447), .O(n10448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__16149.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__16150 (.I0(n8200), .I1(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n10449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16150.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16151 (.I0(n8202), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .O(n10450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16151.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16152 (.I0(n3827), .I1(n8240), .I2(n10400), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n10451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16152.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16153 (.I0(n10449), .I1(n10450), .I2(n10451), .I3(n10436), 
            .O(n10452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__16153.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__16154 (.I0(n10448), .I1(n10441), .I2(n10452), .I3(n10440), 
            .O(n10453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16154.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16155 (.I0(\u_black_pixel_avg/black_pixel_count[25] ), .I1(n8230), 
            .I2(n10089), .O(n10454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16155.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16156 (.I0(n10445), .I1(n10429), .I2(n10453), .I3(n10454), 
            .O(n10455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__16156.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__16210 (.I0(\u_black_pixel_avg/black_pixel_count[30] ), .I1(\u_black_pixel_avg/black_pixel_count[31] ), 
            .O(n10488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16210.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16211 (.I0(\u_black_pixel_avg/black_pixel_count[29] ), .I1(n10488), 
            .O(n10489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16211.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16212 (.I0(n10489), .I1(n9721), .O(n10490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16212.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16680 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[27] ), .I3(\u_black_pixel_avg/black_pixel_count[28] ), 
            .O(n10835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16680.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16681 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n9713), 
            .I2(n10835), .I3(n9722), .O(n10836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__16681.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__16682 (.I0(n9726), .I1(n10836), .O(n10837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16682.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16683 (.I0(\u_black_pixel_avg/black_pixel_count[0] ), .I1(n9744), 
            .I2(n10837), .I3(lcd_vs), .O(n10838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__16683.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__16698 (.I0(\u_black_pixel_avg/y_sum[9] ), .I1(\u_black_pixel_avg/y_sum[8] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16698.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16699 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2862), 
            .I2(\u_black_pixel_avg/y_sum[8] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16699.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16700 (.I0(\u_black_pixel_avg/y_sum[31] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n10854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__16700.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__16701 (.I0(n9710), .I1(n9728), .I2(n10854), .O(n10855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16701.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16702 (.I0(n9726), .I1(n10836), .I2(n10855), .I3(\u_black_pixel_avg/y_sum[31] ), 
            .O(n10856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__16702.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__16703 (.I0(n9710), .I1(n9728), .I2(n10854), .I3(n2367), 
            .O(n10857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__16703.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__16704 (.I0(\u_black_pixel_avg/y_sum[30] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16704.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16705 (.I0(n10857), .I1(n10836), .I2(n10858), .O(n10859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__16705.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__16706 (.I0(\u_black_pixel_avg/y_sum[30] ), .I1(n9702), 
            .O(n10860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16706.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16707 (.I0(n10860), .I1(n9714), .I2(n9709), .O(n10861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__16707.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__16708 (.I0(n10859), .I1(n10856), .I2(n10861), .O(n10862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16708.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16709 (.I0(\u_black_pixel_avg/y_sum[30] ), .I1(n2369), 
            .I2(n10862), .O(n6764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16709.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16710 (.I0(n9709), .I1(n9714), .I2(n10858), .O(n10863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16710.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16711 (.I0(n9726), .I1(n10836), .I2(n10857), .O(n10864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16711.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16712 (.I0(n10860), .I1(n2368), .I2(n9709), .I3(n9714), 
            .O(n10865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__16712.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__16713 (.I0(n10864), .I1(n10856), .I2(n10863), .I3(n10865), 
            .O(n6762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__16713.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__16714 (.I0(\u_black_pixel_avg/y_sum[29] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16714.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16715 (.I0(n9723), .I1(n9726), .I2(n9729), .O(n10867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16715.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16716 (.I0(n6762), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n10866), .I3(n10867), .O(n10868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__16716.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__16717 (.I0(\u_black_pixel_avg/y_sum[29] ), .I1(n9702), 
            .O(n10869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16717.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16718 (.I0(n2372), .I1(n10867), .O(n10870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16718.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16719 (.I0(n6762), .I1(n10869), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n10870), .O(n10871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b00 */ ;
    defparam LUT__16719.LUTMASK = 16'h2b00;
    EFX_LUT4 LUT__16720 (.I0(n10868), .I1(n6764), .I2(n10871), .O(n6769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__16720.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__16721 (.I0(n6764), .I1(n10868), .I2(n10871), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__16721.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__16722 (.I0(\u_black_pixel_avg/y_sum[28] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16722.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16723 (.I0(n10869), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n2369), .O(n10874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__16723.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__16724 (.I0(\u_black_pixel_avg/y_sum[31] ), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[2] ), .I3(\u_black_pixel_avg/y_sum[30] ), 
            .O(n10875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__16724.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__16725 (.I0(n10875), .I1(n10869), .I2(n10866), .O(n10876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__16725.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__16726 (.I0(n10856), .I1(n10859), .I2(n10874), .I3(n10876), 
            .O(n10877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16726.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16727 (.I0(n10877), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n6762), .I3(n10867), .O(n10878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__16727.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__16728 (.I0(\u_black_pixel_avg/y_sum[29] ), .I1(n2374), 
            .I2(n10873), .I3(n10878), .O(n10879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__16728.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__16729 (.I0(\u_black_pixel_avg/y_sum[28] ), .I1(n9702), 
            .O(n10880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16729.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16730 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6762), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n9745), .O(n10881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__16730.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__16731 (.I0(n10872), .I1(n10879), .I2(n10880), .I3(n10881), 
            .O(n10882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__16731.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__16732 (.I0(n9741), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n10877), .I3(n2371), .O(n10883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__16732.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__16733 (.I0(n10867), .I1(n6762), .I2(n2371), .I3(n10883), 
            .O(n6767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc4fc */ ;
    defparam LUT__16733.LUTMASK = 16'hc4fc;
    EFX_LUT4 LUT__16734 (.I0(n10866), .I1(n6762), .I2(n10867), .O(n10884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__16734.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__16735 (.I0(n10884), .I1(n6764), .I2(n10871), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__16735.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__16736 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6767), 
            .I2(n10885), .I3(n10881), .O(n10886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__16736.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__16737 (.I0(n6769), .I1(n2377), .I2(n10882), .I3(n10886), 
            .O(n6776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16737.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16738 (.I0(\u_black_pixel_avg/y_sum[28] ), .I1(n2381), 
            .I2(n10882), .I3(n10886), .O(n6780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16738.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16739 (.I0(\u_black_pixel_avg/y_sum[27] ), .I1(n9702), 
            .O(n10887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16739.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16740 (.I0(\u_black_pixel_avg/y_sum[29] ), .I1(n2374), 
            .I2(n10878), .O(n6771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16740.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16741 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6771), 
            .O(n10888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16741.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16742 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n2379), 
            .O(n10889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16742.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16743 (.I0(n10888), .I1(n10889), .I2(n10882), .I3(n10886), 
            .O(n10890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__16743.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__16744 (.I0(\u_black_pixel_avg/y_sum[27] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16744.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16745 (.I0(n10887), .I1(n6780), .I2(n10891), .I3(n10890), 
            .O(n10892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__16745.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__16746 (.I0(n6771), .I1(n2379), .I2(n10882), .I3(n10886), 
            .O(n6778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16746.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16747 (.I0(n6776), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n6778), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n10893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16747.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16748 (.I0(n6767), .I1(n2376), .I2(n10882), .I3(n10886), 
            .O(n6774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16748.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16749 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6774), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6776), .O(n10894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16749.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16750 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6767), 
            .I2(n9745), .O(n10895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16750.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16751 (.I0(n10892), .I1(n10893), .I2(n10894), .I3(n10895), 
            .O(n10896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16751.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16752 (.I0(n6776), .I1(n2384), .I2(n10896), .O(n6785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16752.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16753 (.I0(n6780), .I1(n2388), .I2(n10896), .O(n6789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16753.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16754 (.I0(\u_black_pixel_avg/y_sum[26] ), .I1(n9702), 
            .O(n10897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16754.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16755 (.I0(\u_black_pixel_avg/y_sum[26] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16755.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16756 (.I0(\u_black_pixel_avg/y_sum[27] ), .I1(n2390), 
            .I2(n10898), .I3(n10896), .O(n10899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__16756.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__16757 (.I0(n10897), .I1(n10899), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n6789), .O(n10900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__16757.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__16758 (.I0(n2386), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n2388), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n10901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16758.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16759 (.I0(n2384), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n10901), .O(n10902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__16759.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__16760 (.I0(n6778), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16760.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16761 (.I0(n6774), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6776), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16761.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16762 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6780), 
            .I2(n10903), .I3(n10904), .O(n10905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__16762.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__16763 (.I0(n10905), .I1(n10902), .I2(n10896), .O(n10906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__16763.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__16764 (.I0(n6774), .I1(n2383), .I2(n10896), .O(n6783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16764.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16765 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6776), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6778), .O(n10907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16765.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16766 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n2384), .I3(n2386), .O(n10908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16766.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16767 (.I0(n10907), .I1(n10904), .I2(n10908), .I3(n10896), 
            .O(n10909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__16767.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__16768 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6783), 
            .I2(n10909), .O(n10910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__16768.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__16769 (.I0(n10906), .I1(n10900), .I2(n10910), .I3(n9775), 
            .O(n10911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__16769.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__16770 (.I0(n6785), .I1(n2393), .I2(n10911), .O(n6796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16770.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16771 (.I0(\u_black_pixel_avg/y_sum[26] ), .I1(n2401), 
            .I2(n10911), .O(n6804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16771.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16772 (.I0(\u_black_pixel_avg/y_sum[25] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16772.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16773 (.I0(\u_black_pixel_avg/y_sum[27] ), .I1(n2390), 
            .I2(n10896), .O(n6791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16773.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16774 (.I0(n6791), .I1(n2399), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n10911), .O(n10913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16774.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16775 (.I0(n6804), .I1(n10912), .I2(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I3(n10913), .O(n10914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__16775.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__16776 (.I0(n6791), .I1(n2399), .I2(n10911), .O(n6802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16776.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16777 (.I0(n6789), .I1(n2397), .I2(n10911), .O(n6800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16777.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16778 (.I0(n6800), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n6802), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n10915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16778.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16779 (.I0(n6778), .I1(n2386), .I2(n10896), .O(n6787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16779.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16780 (.I0(n6787), .I1(n2395), .I2(n10911), .O(n6798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16780.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16781 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6798), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6800), .O(n10916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16781.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16782 (.I0(n6796), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6798), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16782.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16783 (.I0(n10914), .I1(n10915), .I2(n10916), .I3(n10917), 
            .O(n10918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16783.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16784 (.I0(n6783), .I1(n2392), .I2(n10911), .O(n6794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16784.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16785 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6794), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6796), .O(n10919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16785.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16786 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6783), 
            .I2(n9774), .O(n10920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16786.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16787 (.I0(n10919), .I1(n10918), .I2(n10920), .O(n10921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16787.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16788 (.I0(n6796), .I1(n2404), .I2(n10921), .O(n6809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16788.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16789 (.I0(\u_black_pixel_avg/y_sum[24] ), .I1(n9702), 
            .O(n10922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16789.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16790 (.I0(\u_black_pixel_avg/y_sum[25] ), .I1(n2414), 
            .I2(n10922), .I3(n10921), .O(n10923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16790.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16791 (.I0(\u_black_pixel_avg/y_sum[24] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16791.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16792 (.I0(n10924), .I1(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I2(n10920), .I3(\u_black_pixel_avg/y_sum[25] ), .O(n10925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8ee */ ;
    defparam LUT__16792.LUTMASK = 16'he8ee;
    EFX_LUT4 LUT__16793 (.I0(n6804), .I1(n2412), .I2(n10921), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16793.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16794 (.I0(n6802), .I1(n2410), .I2(n10921), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16794.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16795 (.I0(n10925), .I1(n10923), .I2(n10926), .I3(n10927), 
            .O(n10928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16795.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16796 (.I0(n6802), .I1(n2410), .I2(n10921), .O(n6815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16796.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16797 (.I0(n6804), .I1(n2412), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n10921), .O(n10929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16797.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16798 (.I0(n6800), .I1(n2408), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n10921), .O(n10930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16798.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16799 (.I0(n6815), .I1(n10929), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n10930), .O(n10931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__16799.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__16800 (.I0(n6800), .I1(n2408), .I2(n10921), .I3(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n10932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16800.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16801 (.I0(n6798), .I1(n2406), .I2(n10921), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n10933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16801.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16802 (.I0(n2404), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n10934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16802.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16803 (.I0(n6785), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n10935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16803.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16804 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6783), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n9773), .O(n10936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__16804.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__16805 (.I0(n10935), .I1(n10934), .I2(n10921), .I3(n10936), 
            .O(n10937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16805.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16806 (.I0(n10932), .I1(n10933), .I2(n10937), .O(n10938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__16806.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__16807 (.I0(n6796), .I1(n2404), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n10921), .O(n10939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16807.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16808 (.I0(n6798), .I1(n2406), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n10921), .O(n10940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16808.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16809 (.I0(n6794), .I1(n2403), .I2(n10921), .I3(n9774), 
            .O(n10941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__16809.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__16810 (.I0(n10940), .I1(n10939), .I2(n10937), .I3(n10941), 
            .O(n10942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__16810.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__16811 (.I0(n10928), .I1(n10931), .I2(n10938), .I3(n10942), 
            .O(n10943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16811.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16812 (.I0(n2417), .I1(n6809), .I2(n10943), .O(n6824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16812.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16813 (.I0(n6804), .I1(n2412), .I2(n10921), .O(n6817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16813.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16814 (.I0(n2425), .I1(n6817), .I2(n10943), .O(n6832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16814.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16815 (.I0(n2423), .I1(n6815), .I2(n10943), .O(n6830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16815.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16816 (.I0(n6800), .I1(n2408), .I2(n10921), .O(n6813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16816.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16817 (.I0(n2421), .I1(n6813), .I2(n10943), .O(n6828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16817.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16818 (.I0(n6828), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6830), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16818.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16819 (.I0(\u_black_pixel_avg/y_sum[25] ), .I1(n2414), 
            .I2(n10921), .O(n6819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16819.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16820 (.I0(n2427), .I1(n6819), .I2(n10943), .O(n6834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16820.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16821 (.I0(\u_black_pixel_avg/y_sum[23] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__16821.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__16822 (.I0(n2429), .I1(\u_black_pixel_avg/y_sum[24] ), 
            .I2(n10945), .I3(n10943), .O(n10946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16822.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16823 (.I0(\u_black_pixel_avg/y_sum[23] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16823.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16824 (.I0(n6834), .I1(n10946), .I2(n10947), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe */ ;
    defparam LUT__16824.LUTMASK = 16'ha8fe;
    EFX_LUT4 LUT__16825 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6832), 
            .I2(n10944), .I3(n10948), .O(n10949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__16825.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__16826 (.I0(n6830), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n6832), .O(n10950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16826.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16827 (.I0(n10950), .I1(n6828), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n10951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__16827.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__16828 (.I0(n6798), .I1(n2406), .I2(n10921), .O(n6811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16828.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16829 (.I0(n2419), .I1(n6811), .I2(n10943), .O(n6826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16829.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16830 (.I0(n6794), .I1(n2403), .I2(n10921), .O(n6807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16830.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16831 (.I0(n2416), .I1(n6807), .I2(n10943), .O(n6822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16831.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16832 (.I0(n6824), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6822), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16832.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16833 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6826), 
            .I2(n9773), .I3(n10952), .O(n10953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__16833.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__16834 (.I0(n6824), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[6] ), .I3(n6826), .O(n10954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16834.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16835 (.I0(n10954), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n6822), .I3(n9773), .O(n10955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__16835.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__16836 (.I0(n10949), .I1(n10951), .I2(n10953), .I3(n10955), 
            .O(n10956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__16836.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__16837 (.I0(n2432), .I1(n6824), .I2(n10956), .O(n6841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16837.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16838 (.I0(n2440), .I1(n6832), .I2(n10956), .O(n6849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16838.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16839 (.I0(n2442), .I1(n6834), .I2(n10956), .O(n6851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16839.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16840 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6851), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n6849), .O(n10957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16840.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16841 (.I0(n2429), .I1(\u_black_pixel_avg/y_sum[24] ), 
            .I2(n10943), .O(n6836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16841.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16842 (.I0(n2444), .I1(n6836), .I2(n10956), .O(n6853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16842.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16843 (.I0(\u_black_pixel_avg/y_sum[22] ), .I1(n9702), 
            .O(n10958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16843.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16844 (.I0(\u_black_pixel_avg/y_sum[22] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16844.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16845 (.I0(n2446), .I1(\u_black_pixel_avg/y_sum[23] ), 
            .I2(n10959), .I3(n10956), .O(n10960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__16845.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__16846 (.I0(n6853), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n10958), .I3(n10960), .O(n10961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hddd4 */ ;
    defparam LUT__16846.LUTMASK = 16'hddd4;
    EFX_LUT4 LUT__16847 (.I0(n2438), .I1(n6830), .I2(n10956), .O(n6847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16847.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16848 (.I0(n6832), .I1(n6834), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n10962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16848.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16849 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2440), 
            .I2(n2442), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n10963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16849.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16850 (.I0(n10963), .I1(n10962), .I2(n10956), .O(n10964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16850.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16851 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6847), 
            .I2(n10964), .O(n10965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16851.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16852 (.I0(n10961), .I1(n10957), .I2(n10965), .O(n10966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__16852.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__16853 (.I0(n2436), .I1(n6828), .I2(n10956), .O(n6845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16853.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16854 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6845), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6847), .O(n10967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16854.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16855 (.I0(n2434), .I1(n6826), .I2(n10956), .O(n6843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16855.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16856 (.I0(n2432), .I1(n6824), .I2(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I3(n10956), .O(n10968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16856.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16857 (.I0(n2431), .I1(n6822), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(n10956), .O(n10969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16857.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16858 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6843), 
            .I2(n10968), .I3(n10969), .O(n10970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__16858.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__16859 (.I0(n6845), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n6843), .I3(\u_black_pixel_avg/black_pixel_count[7] ), .O(n10971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16859.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16860 (.I0(n2431), .I1(n6822), .I2(n10956), .O(n6839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16860.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16861 (.I0(n6839), .I1(n6841), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16861.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16862 (.I0(n10971), .I1(n10970), .I2(n10972), .I3(n9838), 
            .O(n10973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__16862.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__16863 (.I0(n10966), .I1(n10970), .I2(n10967), .I3(n10973), 
            .O(n10974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__16863.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__16864 (.I0(n6841), .I1(n2449), .I2(n10974), .O(n6860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16864.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16865 (.I0(n2446), .I1(\u_black_pixel_avg/y_sum[23] ), 
            .I2(n10956), .O(n6855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16865.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16866 (.I0(n6855), .I1(n2463), .I2(n10974), .O(n6874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16866.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16867 (.I0(\u_black_pixel_avg/y_sum[22] ), .I1(n2465), 
            .I2(n10974), .O(n6876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16867.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16868 (.I0(n6876), .I1(\u_black_pixel_avg/y_sum[21] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n10975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16868.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16869 (.I0(n6855), .I1(n2463), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n10974), .O(n10976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16869.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16870 (.I0(n6851), .I1(n2459), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n10974), .O(n10977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16870.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16871 (.I0(n6853), .I1(n2461), .I2(n10974), .O(n6872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16871.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16872 (.I0(n6872), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n10977), .I3(n10976), .O(n10978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16872.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16873 (.I0(n6874), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n10975), .I3(n10978), .O(n10979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16873.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16874 (.I0(n2459), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n2461), .I3(n10974), .O(n10980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d33 */ ;
    defparam LUT__16874.LUTMASK = 16'h0d33;
    EFX_LUT4 LUT__16875 (.I0(n6851), .I1(n10980), .I2(n6853), .I3(n10974), 
            .O(n10981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcc07 */ ;
    defparam LUT__16875.LUTMASK = 16'hcc07;
    EFX_LUT4 LUT__16876 (.I0(n6851), .I1(n2459), .I2(n10974), .O(n6870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16876.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16877 (.I0(n6849), .I1(n2457), .I2(n10974), .O(n6868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16877.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16878 (.I0(n6868), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6870), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n10982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16878.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16879 (.I0(n6847), .I1(n2455), .I2(n10974), .O(n6866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16879.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16880 (.I0(n6845), .I1(n2453), .I2(n10974), .O(n6864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16880.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16881 (.I0(n6864), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n6866), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n10983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16881.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16882 (.I0(n10981), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n10982), .I3(n10983), .O(n10984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__16882.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__16883 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6868), 
            .I2(\u_black_pixel_avg/black_pixel_count[6] ), .I3(n6866), .O(n10985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16883.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16884 (.I0(n6839), .I1(n2448), .I2(n10974), .O(n6858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16884.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16885 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6858), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6860), .O(n10986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16885.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16886 (.I0(n6843), .I1(n2451), .I2(n10974), .O(n6862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16886.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16887 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6862), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6864), .O(n10987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16887.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16888 (.I0(n10985), .I1(n10983), .I2(n10986), .I3(n10987), 
            .O(n10988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__16888.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__16889 (.I0(n6860), .I1(n6862), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n10989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16889.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16890 (.I0(n10989), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n6858), .I3(n9837), .O(n10990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__16890.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__16891 (.I0(n10979), .I1(n10984), .I2(n10988), .I3(n10990), 
            .O(n10991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__16891.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__16892 (.I0(n6860), .I1(n2468), .I2(n10991), .O(n6881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16892.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16893 (.I0(n6872), .I1(n2480), .I2(n10991), .O(n6893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16893.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16894 (.I0(n6874), .I1(n2482), .I2(n10991), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n10992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16894.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16895 (.I0(n6870), .I1(n2478), .I2(n10991), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n10993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16895.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16896 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6893), 
            .I2(n10992), .I3(n10993), .O(n10994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16896.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16897 (.I0(n6876), .I1(n2484), .I2(n10991), .O(n6897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16897.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16898 (.I0(\u_black_pixel_avg/y_sum[20] ), .I1(n9702), 
            .O(n10995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16898.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16899 (.I0(\u_black_pixel_avg/y_sum[21] ), .I1(n2486), 
            .I2(n10995), .I3(n10991), .O(n10996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16899.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16900 (.I0(\u_black_pixel_avg/y_sum[20] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n10997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__16900.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__16901 (.I0(n6897), .I1(n10996), .I2(n10997), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n10998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe */ ;
    defparam LUT__16901.LUTMASK = 16'ha8fe;
    EFX_LUT4 LUT__16902 (.I0(n6874), .I1(n2482), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n10991), .O(n10999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16902.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16903 (.I0(n6893), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n10999), .I3(n10993), .O(n11000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__16903.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__16904 (.I0(n6870), .I1(n2478), .I2(n10991), .O(n6891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16904.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16905 (.I0(n6868), .I1(n2476), .I2(n10991), .O(n6889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16905.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16906 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6889), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n6891), .O(n11001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16906.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16907 (.I0(n10998), .I1(n10994), .I2(n11000), .I3(n11001), 
            .O(n11002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__16907.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__16908 (.I0(n6862), .I1(n2470), .I2(n10991), .O(n6883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16908.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16909 (.I0(n6883), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16909.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16910 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6858), 
            .I2(n9875), .O(n11004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16910.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16911 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6881), 
            .I2(n11004), .O(n11005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16911.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16912 (.I0(n6866), .I1(n2474), .I2(n10991), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16912.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16913 (.I0(n6864), .I1(n2472), .I2(n10991), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n11007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16913.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16914 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6889), 
            .I2(n11006), .I3(n11007), .O(n11008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16914.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16915 (.I0(n11003), .I1(n11005), .I2(n11008), .O(n11009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__16915.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__16916 (.I0(n6864), .I1(n2472), .I2(n10991), .O(n6885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16916.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16917 (.I0(n6866), .I1(n2474), .I2(n10991), .O(n6887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16917.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16918 (.I0(n6885), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n6887), .O(n11010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16918.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16919 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6883), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n6881), 
            .O(n11011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16919.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16920 (.I0(n11003), .I1(n11010), .I2(n11011), .I3(n11005), 
            .O(n11012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__16920.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__16921 (.I0(n6858), .I1(n2467), .I2(n10991), .O(n6879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16921.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16922 (.I0(n6879), .I1(n9837), .O(n11013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16922.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16923 (.I0(n11009), .I1(n11002), .I2(n11012), .I3(n11013), 
            .O(n11014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16923.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16924 (.I0(n2489), .I1(n6881), .I2(n11014), .O(n6904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16924.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16925 (.I0(n2495), .I1(n6887), .I2(n11014), .O(n6910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16925.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16926 (.I0(n2497), .I1(n6889), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11014), .O(n11015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16926.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16927 (.I0(n2493), .I1(n6885), .I2(n11014), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16927.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16928 (.I0(n6910), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n11015), .I3(n11016), .O(n11017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__16928.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__16929 (.I0(n2493), .I1(n6885), .I2(n11014), .O(n6908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16929.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16930 (.I0(n2491), .I1(n6883), .I2(n11014), .O(n6906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16930.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16931 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6906), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n6908), .O(n11018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16931.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16932 (.I0(n11009), .I1(n11002), .I2(n11012), .I3(n9837), 
            .O(n11019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16932.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16933 (.I0(n11009), .I1(n11002), .I2(n11012), .I3(n6879), 
            .O(n11020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__16933.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__16934 (.I0(n2488), .I1(n11019), .I2(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I3(n11020), .O(n11021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__16934.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__16935 (.I0(n2489), .I1(n6881), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(n11014), .O(n11022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16935.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16936 (.I0(n11021), .I1(n11022), .O(n11023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16936.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16937 (.I0(n6883), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n6881), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16937.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16938 (.I0(n2489), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n2491), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16938.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16939 (.I0(n11025), .I1(n11024), .I2(n11014), .O(n11026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__16939.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__16940 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6879), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n9744), 
            .O(n11027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__16940.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__16941 (.I0(n11021), .I1(n11022), .I2(n11026), .I3(n11027), 
            .O(n11028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__16941.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__16942 (.I0(n11017), .I1(n11023), .I2(n11018), .I3(n11028), 
            .O(n11029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__16942.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__16943 (.I0(n2505), .I1(n6897), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n11014), .O(n11030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16943.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16944 (.I0(n6874), .I1(n2482), .I2(n10991), .O(n6895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16944.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16945 (.I0(n2503), .I1(n6895), .I2(n11014), .O(n6918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16945.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16946 (.I0(n2501), .I1(n6893), .I2(n11014), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n11031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16946.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16947 (.I0(n11030), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n6918), .I3(n11031), .O(n11032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__16947.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__16948 (.I0(n2499), .I1(n6891), .I2(n11014), .O(n6914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16948.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16949 (.I0(n2501), .I1(n6893), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n11014), .O(n11033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16949.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16950 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2509), 
            .I2(\u_black_pixel_avg/y_sum[19] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__16950.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__16951 (.I0(n2501), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n11035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16951.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16952 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n2507), 
            .I2(n11034), .I3(n11035), .O(n11036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__16952.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__16953 (.I0(n2503), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n2505), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n11037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16953.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16954 (.I0(\u_black_pixel_avg/y_sum[21] ), .I1(n2486), 
            .I2(n10991), .O(n6899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16954.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16955 (.I0(\u_black_pixel_avg/y_sum[20] ), .I1(\u_black_pixel_avg/y_sum[19] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__16955.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__16956 (.I0(n6893), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n6897), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n11039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16956.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16957 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6895), 
            .I2(n11039), .O(n11040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__16957.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__16958 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6899), 
            .I2(n11038), .I3(n11040), .O(n11041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd400 */ ;
    defparam LUT__16958.LUTMASK = 16'hd400;
    EFX_LUT4 LUT__16959 (.I0(n11037), .I1(n11036), .I2(n11041), .I3(n11014), 
            .O(n11042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__16959.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__16960 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6914), 
            .I2(n11033), .I3(n11042), .O(n11043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__16960.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__16961 (.I0(n2495), .I1(n6887), .I2(n11014), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n11044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16961.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16962 (.I0(n2499), .I1(n6891), .I2(n11014), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16962.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16963 (.I0(n2497), .I1(n6889), .I2(n11014), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16963.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16964 (.I0(n11016), .I1(n11044), .I2(n11045), .I3(n11046), 
            .O(n11047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16964.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16965 (.I0(n11043), .I1(n11032), .I2(n11028), .I3(n11047), 
            .O(n11048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__16965.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__16966 (.I0(n11029), .I1(n11048), .O(n11049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16966.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16967 (.I0(n2512), .I1(n6904), .I2(n11049), .O(n6929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16967.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16968 (.I0(n6908), .I1(n2516), .I2(n11029), .I3(n11048), 
            .O(n6933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16968.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16969 (.I0(n6910), .I1(n2518), .I2(n11029), .I3(n11048), 
            .O(n6935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16969.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16970 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6935), 
            .O(n11050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16970.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16971 (.I0(n6906), .I1(n2514), .I2(n11029), .I3(n11048), 
            .O(n6931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16971.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16972 (.I0(n6933), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n6931), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16972.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16973 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n6933), 
            .I2(n11050), .I3(n11051), .O(n11052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__16973.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__16974 (.I0(n2522), .I1(n6914), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11049), .O(n11053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16974.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16975 (.I0(n2497), .I1(n6889), .I2(n11014), .O(n6912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16975.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16976 (.I0(n6912), .I1(n2520), .I2(n11029), .I3(n11048), 
            .O(n6937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__16976.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__16977 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6937), 
            .O(n11054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16977.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16978 (.I0(n6937), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n6935), .I3(\u_black_pixel_avg/black_pixel_count[9] ), .O(n11055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16978.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16979 (.I0(n11054), .I1(n11053), .I2(n11051), .I3(n11055), 
            .O(n11056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__16979.LUTMASK = 16'he000;
    EFX_LUT4 LUT__16980 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6931), 
            .O(n11057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16980.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16981 (.I0(n2488), .I1(n11019), .I2(n11020), .O(n6902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__16981.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__16982 (.I0(n2511), .I1(n6902), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n11049), .O(n11058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16982.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16983 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6929), 
            .I2(n11057), .I3(n11058), .O(n11059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__16983.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__16984 (.I0(n2511), .I1(n6902), .I2(n11049), .O(n6927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16984.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16985 (.I0(n2512), .I1(n6904), .I2(n11049), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__16985.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__16986 (.I0(n6927), .I1(n11060), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n9744), .O(n11061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b00 */ ;
    defparam LUT__16986.LUTMASK = 16'h2b00;
    EFX_LUT4 LUT__16987 (.I0(n11056), .I1(n11052), .I2(n11059), .I3(n11061), 
            .O(n11062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__16987.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__16988 (.I0(n2509), .I1(\u_black_pixel_avg/y_sum[20] ), 
            .I2(n11014), .O(n6924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16988.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16989 (.I0(n2532), .I1(n6924), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n11049), .O(n11063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16989.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16990 (.I0(\u_black_pixel_avg/y_sum[18] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/y_sum[19] ), 
            .O(n11064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__16990.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__16991 (.I0(\u_black_pixel_avg/y_sum[18] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(n2534), .O(n11065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__16991.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__16992 (.I0(\u_black_pixel_avg/y_sum[18] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__16992.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__16993 (.I0(n11065), .I1(n11064), .I2(n11066), .I3(n11049), 
            .O(n11067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__16993.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__16994 (.I0(n6918), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n11068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16994.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16995 (.I0(n2505), .I1(n6897), .I2(n11014), .O(n6920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16995.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16996 (.I0(n6924), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n6920), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16996.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16997 (.I0(n2526), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2532), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n11070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__16997.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__16998 (.I0(n2528), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n11070), .O(n11071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__16998.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__16999 (.I0(n11068), .I1(n11069), .I2(n11071), .I3(n11049), 
            .O(n11072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__16999.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__17000 (.I0(n2507), .I1(n6899), .I2(n11014), .O(n6922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17000.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17001 (.I0(n6922), .I1(n2530), .I2(n11029), .I3(n11048), 
            .O(n6947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17001.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17002 (.I0(n6947), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n11073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17002.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17003 (.I0(n11067), .I1(n11063), .I2(n11072), .I3(n11073), 
            .O(n11074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__17003.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__17004 (.I0(n11068), .I1(n6920), .O(n11075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17004.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17005 (.I0(n2526), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2528), .O(n11076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17005.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17006 (.I0(n11075), .I1(n11076), .I2(n11029), .I3(n11048), 
            .O(n11077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17006.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17007 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6947), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n11077), 
            .O(n11078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__17007.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__17008 (.I0(n11068), .I1(n6922), .O(n11079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17008.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17009 (.I0(n2526), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2530), .O(n11080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17009.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17010 (.I0(n11080), .I1(n11079), .I2(n11049), .I3(n9727), 
            .O(n11081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__17010.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__17011 (.I0(n2526), .I1(n6918), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n11049), .O(n11082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17011.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17012 (.I0(n2501), .I1(n6893), .I2(n11014), .O(n6916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17012.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17013 (.I0(n2524), .I1(n6916), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n11049), .O(n11083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17013.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17014 (.I0(n11078), .I1(n11081), .I2(n11082), .I3(n11083), 
            .O(n11084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17014.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17015 (.I0(n2524), .I1(n6916), .I2(n11049), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17015.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17016 (.I0(n2522), .I1(n6914), .I2(n11049), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17016.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17017 (.I0(n11085), .I1(n11086), .I2(n11051), .I3(n11055), 
            .O(n11087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__17017.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__17018 (.I0(n11084), .I1(n11074), .I2(n11061), .I3(n11087), 
            .O(n11088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__17018.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__17019 (.I0(n11062), .I1(n11088), .O(n11089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__17019.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__17020 (.I0(n2537), .I1(n6929), .I2(n11089), .O(n6956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17020.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17021 (.I0(n2553), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2555), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17021.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17022 (.I0(n2557), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n2559), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n11091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17022.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17023 (.I0(n2534), .I1(\u_black_pixel_avg/y_sum[19] ), 
            .I2(n11049), .O(n6951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17023.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17024 (.I0(n2532), .I1(n6924), .I2(n11049), .O(n6949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17024.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17025 (.I0(n6949), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n6951), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n11092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17025.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17026 (.I0(n2528), .I1(n6920), .I2(n11049), .O(n6945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17026.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17027 (.I0(n6947), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n6945), .I3(\u_black_pixel_avg/black_pixel_count[5] ), .O(n11093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17027.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17028 (.I0(n11092), .I1(n11093), .O(n11094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17028.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17029 (.I0(n11091), .I1(n11090), .I2(n11094), .I3(n11089), 
            .O(n11095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__17029.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__17030 (.I0(n6951), .I1(n2559), .I2(n11062), .I3(n11088), 
            .O(n6978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17030.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17031 (.I0(\u_black_pixel_avg/y_sum[17] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17031.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17032 (.I0(\u_black_pixel_avg/y_sum[17] ), .I1(n9702), 
            .I2(\u_black_pixel_avg/y_sum[18] ), .O(n11097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17032.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17033 (.I0(\u_black_pixel_avg/y_sum[17] ), .I1(n9702), 
            .I2(n2561), .O(n11098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17033.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17034 (.I0(n11097), .I1(n11098), .I2(n11062), .I3(n11088), 
            .O(n11099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17034.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17035 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6978), 
            .I2(n11096), .I3(n11099), .O(n11100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__17035.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__17036 (.I0(n2553), .I1(n6945), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n11089), .O(n11101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17036.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17037 (.I0(n2526), .I1(n6918), .I2(n11049), .O(n6943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17037.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17038 (.I0(n6943), .I1(n2551), .I2(n11062), .I3(n11088), 
            .O(n6970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17038.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17039 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2555), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n2557), .O(n11102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17039.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17040 (.I0(n11088), .I1(n11062), .I2(n11102), .I3(n11090), 
            .O(n11103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__17040.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__17041 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n6947), 
            .O(n11104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17041.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17042 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n6949), 
            .I2(n11104), .I3(n11093), .O(n11105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__17042.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__17043 (.I0(n11062), .I1(n11088), .I2(n11105), .O(n11106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17043.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17044 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6970), 
            .I2(n11103), .I3(n11106), .O(n11107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__17044.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__17045 (.I0(n11100), .I1(n11095), .I2(n11101), .I3(n11107), 
            .O(n11108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__17045.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__17046 (.I0(n2524), .I1(n6916), .I2(n11049), .O(n6941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17046.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17047 (.I0(n6941), .I1(n2549), .I2(n11062), .I3(n11088), 
            .O(n6968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17047.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17048 (.I0(n6970), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17048.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17049 (.I0(n6933), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17049.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17050 (.I0(n2541), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17050.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17051 (.I0(n11110), .I1(n11111), .I2(n11062), .I3(n11088), 
            .O(n11112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17051.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17052 (.I0(n6935), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17052.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17053 (.I0(n2543), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17053.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17054 (.I0(n11113), .I1(n11114), .I2(n11062), .I3(n11088), 
            .O(n11115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17054.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17055 (.I0(n2522), .I1(n6914), .I2(n11049), .O(n6939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17055.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17056 (.I0(n6939), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n11116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17056.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17057 (.I0(n2547), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n11117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17057.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17058 (.I0(n11116), .I1(n11117), .I2(n11062), .I3(n11088), 
            .O(n11118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17058.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17059 (.I0(n6937), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17059.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17060 (.I0(n2545), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17060.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17061 (.I0(n11119), .I1(n11120), .I2(n11062), .I3(n11088), 
            .O(n11121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17061.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17062 (.I0(n11112), .I1(n11115), .I2(n11118), .I3(n11121), 
            .O(n11122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__17062.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__17063 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6968), 
            .I2(n11109), .I3(n11122), .O(n11123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17063.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17064 (.I0(n2543), .I1(n6935), .I2(n11089), .O(n6962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17064.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17065 (.I0(n2545), .I1(n6937), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(n11089), .O(n11124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17065.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17066 (.I0(n6962), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n11124), .I3(n11112), .O(n11125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__17066.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__17067 (.I0(n6939), .I1(n2547), .I2(n11062), .I3(n11088), 
            .O(n6966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17067.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17068 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6968), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n6966), .O(n11126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17068.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17069 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n6929), 
            .O(n11127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17069.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17070 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n2537), 
            .O(n11128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17070.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17071 (.I0(n6927), .I1(n9744), .O(n11129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17071.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17072 (.I0(n11129), .I1(n2536), .I2(n11062), .I3(n11088), 
            .O(n11130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17072.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17073 (.I0(n11128), .I1(n11127), .I2(n11130), .I3(n11089), 
            .O(n11131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17073.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17074 (.I0(n6933), .I1(n2541), .I2(n11062), .I3(n11088), 
            .O(n6960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17074.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17075 (.I0(n6931), .I1(n2539), .I2(n11062), .I3(n11088), 
            .O(n6958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17075.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17076 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6958), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n6960), 
            .O(n11132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17076.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17077 (.I0(n11126), .I1(n11122), .I2(n11131), .I3(n11132), 
            .O(n11133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__17077.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__17078 (.I0(n11123), .I1(n11108), .I2(n11125), .I3(n11133), 
            .O(n11134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17078.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17079 (.I0(n6958), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17079.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17080 (.I0(n2536), .I1(n6927), .I2(n11089), .O(n6954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17080.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17081 (.I0(n6954), .I1(n6956), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[13] ), .O(n11136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17081.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17082 (.I0(n11135), .I1(n11131), .I2(n11136), .I3(n9978), 
            .O(n11137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__17082.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__17083 (.I0(n11134), .I1(n11137), .O(n11138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17083.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17084 (.I0(n6956), .I1(n2564), .I2(n11138), .O(n6985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17084.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17085 (.I0(n2590), .I1(\u_black_pixel_avg/y_sum[17] ), 
            .I2(n11134), .I3(n11137), .O(n7011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17085.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17086 (.I0(\u_black_pixel_avg/y_sum[16] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17086.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17087 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n2588), 
            .O(n11140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17087.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17088 (.I0(n2561), .I1(\u_black_pixel_avg/y_sum[18] ), 
            .I2(n11089), .O(n6980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17088.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17089 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n6980), 
            .O(n11141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17089.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17090 (.I0(n11140), .I1(n11141), .I2(n11134), .I3(n11137), 
            .O(n11142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17090.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17091 (.I0(n7011), .I1(n11139), .I2(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I3(n11142), .O(n11143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd400 */ ;
    defparam LUT__17091.LUTMASK = 16'hd400;
    EFX_LUT4 LUT__17092 (.I0(n2588), .I1(n6980), .I2(n11134), .I3(n11137), 
            .O(n7009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17092.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17093 (.I0(n2586), .I1(n6978), .I2(n11134), .I3(n11137), 
            .O(n7007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17093.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17094 (.I0(n7007), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n7009), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n11144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17094.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17095 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n2578), 
            .O(n11145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17095.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17096 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n6970), 
            .O(n11146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17096.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17097 (.I0(n11145), .I1(n11146), .I2(n11134), .I3(n11137), 
            .O(n11147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17097.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17098 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n2576), 
            .O(n11148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17098.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17099 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6968), 
            .O(n11149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17099.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17100 (.I0(n11148), .I1(n11149), .I2(n11134), .I3(n11137), 
            .O(n11150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17100.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17101 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n7007), 
            .I2(n11147), .I3(n11150), .O(n11151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__17101.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__17102 (.I0(n2557), .I1(n6949), .I2(n11089), .O(n6976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17102.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17103 (.I0(n2584), .I1(n6976), .I2(n11134), .I3(n11137), 
            .O(n7005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17103.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17104 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n2580), 
            .O(n11152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17104.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17105 (.I0(n2553), .I1(n6945), .I2(n11089), .O(n6972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17105.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17106 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n6972), 
            .O(n11153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17106.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17107 (.I0(n11152), .I1(n11153), .I2(n11134), .I3(n11137), 
            .O(n11154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17107.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17108 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n2582), 
            .O(n11155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17108.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17109 (.I0(n2555), .I1(n6947), .I2(n11089), .O(n6974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17109.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17110 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n6974), 
            .O(n11156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17110.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17111 (.I0(n11155), .I1(n11156), .I2(n11134), .I3(n11137), 
            .O(n11157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17111.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17112 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7005), 
            .I2(n11154), .I3(n11157), .O(n11158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__17112.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__17113 (.I0(n11144), .I1(n11143), .I2(n11151), .I3(n11158), 
            .O(n11159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__17113.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__17114 (.I0(n2582), .I1(n6974), .I2(n11134), .I3(n11137), 
            .O(n7003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17114.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17115 (.I0(n7003), .I1(n7005), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17115.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17116 (.I0(n2580), .I1(n6972), .I2(n11134), .I3(n11137), 
            .O(n7001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17116.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17117 (.I0(n2578), .I1(n6970), .I2(n11134), .I3(n11137), 
            .O(n6999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17117.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17118 (.I0(n6999), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n7001), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n11161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17118.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17119 (.I0(n11150), .I1(n11147), .O(n11162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17119.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17120 (.I0(n11160), .I1(n11154), .I2(n11161), .I3(n11162), 
            .O(n11163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17120.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17121 (.I0(n6956), .I1(n2564), .I2(n11138), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17121.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17122 (.I0(n6954), .I1(n2563), .I2(n11138), .O(n6983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17122.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17123 (.I0(n11164), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n6983), .I3(n9977), .O(n11165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__17123.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__17124 (.I0(n2570), .I1(n6962), .I2(n11134), .I3(n11137), 
            .O(n6991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17124.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17125 (.I0(n6991), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17125.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17126 (.I0(n6966), .I1(n2574), .I2(n11138), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17126.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17127 (.I0(n2568), .I1(n6960), .I2(n11134), .I3(n11137), 
            .O(n6989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17127.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17128 (.I0(n2566), .I1(n6958), .I2(n11134), .I3(n11137), 
            .O(n6987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17128.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17129 (.I0(n6987), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n6989), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17129.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17130 (.I0(n2545), .I1(n6937), .I2(n11089), .O(n6964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17130.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17131 (.I0(n2572), .I1(n6964), .I2(n11134), .I3(n11137), 
            .O(n6993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17131.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17132 (.I0(n2576), .I1(n6968), .I2(n11134), .I3(n11137), 
            .O(n6997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17132.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17133 (.I0(n6997), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n6993), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17133.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17134 (.I0(n11166), .I1(n11167), .I2(n11168), .I3(n11169), 
            .O(n11170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__17134.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__17135 (.I0(n11159), .I1(n11163), .I2(n11165), .I3(n11170), 
            .O(n11171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__17135.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__17136 (.I0(n6966), .I1(n2574), .I2(n11138), .I3(n9725), 
            .O(n11172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__17136.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__17137 (.I0(n2574), .I1(n6966), .I2(n11134), .I3(n11137), 
            .O(n11173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17137.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17138 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n11173), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n6993), 
            .O(n11174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__17138.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__17139 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6991), 
            .I2(\u_black_pixel_avg/black_pixel_count[12] ), .I3(n6989), 
            .O(n11175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17139.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17140 (.I0(n11174), .I1(n11172), .I2(n11166), .I3(n11175), 
            .O(n11176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__17140.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__17141 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n6987), 
            .O(n11177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17141.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17142 (.I0(n6954), .I1(n2563), .I2(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I3(n11138), .O(n11178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17142.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17143 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n6985), 
            .I2(n11177), .I3(n11178), .O(n11179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__17143.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__17144 (.I0(n11176), .I1(n11168), .I2(n11179), .I3(n11165), 
            .O(n11180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17144.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17145 (.I0(n11171), .I1(n11180), .O(n11181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__17145.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__17146 (.I0(n2593), .I1(n6985), .I2(n11181), .O(n7016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17146.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17147 (.I0(\u_black_pixel_avg/y_sum[16] ), .I1(n2621), 
            .I2(n11171), .I3(n11180), .O(n7044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17147.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17148 (.I0(\u_black_pixel_avg/y_sum[15] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17148.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17149 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n7011), 
            .O(n11183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17149.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17150 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n2619), 
            .O(n11184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17150.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17151 (.I0(n11183), .I1(n11184), .I2(n11171), .I3(n11180), 
            .O(n11185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17151.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17152 (.I0(n7044), .I1(n11182), .I2(\u_black_pixel_avg/black_pixel_count[1] ), 
            .I3(n11185), .O(n11186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd400 */ ;
    defparam LUT__17152.LUTMASK = 16'hd400;
    EFX_LUT4 LUT__17153 (.I0(n7011), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n7009), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n11187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17153.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17154 (.I0(n2617), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n2619), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n11188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17154.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17155 (.I0(n7005), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n7007), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17155.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17156 (.I0(n2613), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2615), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17156.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17157 (.I0(n11189), .I1(n11190), .I2(n11171), .I3(n11180), 
            .O(n11191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17157.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17158 (.I0(n11188), .I1(n11187), .I2(n11191), .I3(n11181), 
            .O(n11192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17158.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17159 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7007), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n7009), .O(n11193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17159.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17160 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2615), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n2617), .O(n11194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17160.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17161 (.I0(n11194), .I1(n11193), .I2(n11191), .I3(n11181), 
            .O(n11195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17161.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17162 (.I0(n7003), .I1(n2611), .I2(n11171), .I3(n11180), 
            .O(n7034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17162.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17163 (.I0(n7005), .I1(n2613), .I2(n11171), .I3(n11180), 
            .O(n7036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17163.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17164 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n7036), 
            .I2(\u_black_pixel_avg/black_pixel_count[6] ), .I3(n7034), .O(n11196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17164.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17165 (.I0(n11192), .I1(n11186), .I2(n11195), .I3(n11196), 
            .O(n11197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17165.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17166 (.I0(n2609), .I1(n7001), .I2(n11181), .O(n7032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17166.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17167 (.I0(n7034), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17167.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17168 (.I0(n6999), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n6997), .I3(\u_black_pixel_avg/black_pixel_count[9] ), .O(n11199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17168.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17169 (.I0(n2605), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n2607), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17169.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17170 (.I0(n6966), .I1(n2574), .I2(n11138), .O(n6995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17170.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17171 (.I0(n6993), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n6995), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17171.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17172 (.I0(n2601), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n2603), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17172.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17173 (.I0(n11201), .I1(n11202), .I2(n11171), .I3(n11180), 
            .O(n11203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17173.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17174 (.I0(n11200), .I1(n11199), .I2(n11203), .I3(n11181), 
            .O(n11204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17174.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17175 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n7032), 
            .I2(n11198), .I3(n11204), .O(n11205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17175.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17176 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n6999), 
            .O(n11206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17176.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17177 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n7001), 
            .O(n11207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17177.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17178 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n2607), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n2609), .O(n11208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17178.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17179 (.I0(n11207), .I1(n11206), .I2(n11208), .I3(n11181), 
            .O(n11209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__17179.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__17180 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n6997), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n6995), 
            .O(n11210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17180.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17181 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n2603), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n2605), .O(n11211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17181.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17182 (.I0(n11211), .I1(n11210), .I2(n11203), .I3(n11181), 
            .O(n11212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17182.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17183 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n6983), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n6985), 
            .O(n11213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17183.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17184 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n6987), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n6989), 
            .O(n11214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17184.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17185 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n6991), 
            .I2(n11213), .I3(n11214), .O(n11215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__17185.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__17186 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n2592), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n2593), 
            .O(n11216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17186.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17187 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n2595), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n2597), 
            .O(n11217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17187.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17188 (.I0(n2599), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n11216), .I3(n11217), .O(n11218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__17188.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__17189 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n6993), 
            .O(n11219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17189.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17190 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n2601), 
            .O(n11220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17190.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17191 (.I0(n11219), .I1(n11220), .I2(n11171), .I3(n11180), 
            .O(n11221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17191.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17192 (.I0(n11218), .I1(n11215), .I2(n11181), .I3(n11221), 
            .O(n11222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__17192.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__17193 (.I0(n11209), .I1(n11204), .I2(n11212), .I3(n11222), 
            .O(n11223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__17193.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__17194 (.I0(n2597), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n2599), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17194.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17195 (.I0(n2593), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n2595), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17195.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17196 (.I0(n11224), .I1(n11217), .I2(n11225), .I3(n11216), 
            .O(n11226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17196.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17197 (.I0(n6991), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n6989), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n11227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17197.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17198 (.I0(n6987), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n6985), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n11228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17198.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17199 (.I0(n11227), .I1(n11214), .I2(n11228), .I3(n11213), 
            .O(n11229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17199.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17200 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n6983), 
            .I2(n11229), .I3(n9976), .O(n11230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17200.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17201 (.I0(n11226), .I1(n11181), .I2(n11230), .O(n11231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17201.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17202 (.I0(n11197), .I1(n11205), .I2(n11223), .I3(n11231), 
            .O(n11232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17202.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17203 (.I0(n7016), .I1(n2624), .I2(n11232), .O(n7833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17203.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17204 (.I0(n2619), .I1(n7011), .I2(n11181), .O(n7042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17204.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17205 (.I0(n7042), .I1(n2650), .I2(n11232), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n11233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17205.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17206 (.I0(n7044), .I1(n2652), .I2(n11232), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n11234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17206.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17207 (.I0(\u_black_pixel_avg/y_sum[14] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17207.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17208 (.I0(\u_black_pixel_avg/y_sum[15] ), .I1(n2654), 
            .I2(n11235), .I3(n11232), .O(n11236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17208.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17209 (.I0(\u_black_pixel_avg/y_sum[14] ), .I1(n9702), 
            .O(n11237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17209.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17210 (.I0(n11233), .I1(n11234), .I2(n11236), .I3(n11237), 
            .O(n11238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17210.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17211 (.I0(n7042), .I1(n2650), .I2(n11232), .O(n7071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17211.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17212 (.I0(n7044), .I1(n2652), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n11232), .O(n11239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17212.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17213 (.I0(n2617), .I1(n7009), .I2(n11181), .O(n7040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17213.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17214 (.I0(n7040), .I1(n2648), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n11232), .O(n11240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17214.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17215 (.I0(n7071), .I1(n11239), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n11240), .O(n11241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__17215.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__17216 (.I0(n2607), .I1(n6999), .I2(n11181), .O(n7030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17216.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17217 (.I0(n7030), .I1(n2638), .I2(n11232), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17217.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17218 (.I0(n7032), .I1(n2640), .I2(n11232), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n11243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17218.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17219 (.I0(n7036), .I1(n2644), .I2(n11232), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17219.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17220 (.I0(n7034), .I1(n2642), .I2(n11232), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17220.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17221 (.I0(n11242), .I1(n11243), .I2(n11244), .I3(n11245), 
            .O(n11246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17221.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17222 (.I0(n7040), .I1(n2648), .I2(n11232), .O(n7069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17222.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17223 (.I0(n2615), .I1(n7007), .I2(n11181), .O(n7038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17223.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17224 (.I0(n7038), .I1(n2646), .I2(n11232), .O(n7067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17224.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17225 (.I0(n7067), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n7069), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17225.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17226 (.I0(n11241), .I1(n11238), .I2(n11246), .I3(n11247), 
            .O(n11248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__17226.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__17227 (.I0(n7036), .I1(n2644), .I2(n11232), .O(n7065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17227.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17228 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n7067), 
            .I2(\u_black_pixel_avg/black_pixel_count[6] ), .I3(n7065), .O(n11249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17228.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17229 (.I0(n7032), .I1(n2640), .I2(n11232), .O(n7061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17229.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17230 (.I0(n7034), .I1(n2642), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11232), .O(n11250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17230.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17231 (.I0(n7061), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n11250), .I3(n11242), .O(n11251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17231.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17232 (.I0(n7030), .I1(n2638), .I2(n11232), .O(n7059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17232.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17233 (.I0(n2605), .I1(n6997), .I2(n11181), .O(n7028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17233.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17234 (.I0(n7028), .I1(n2636), .I2(n11232), .O(n7057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17234.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17235 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7057), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7059), .O(n11252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17235.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17236 (.I0(n11249), .I1(n11246), .I2(n11251), .I3(n11252), 
            .O(n11253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__17236.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__17237 (.I0(n2599), .I1(n6991), .I2(n11181), .O(n7022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17237.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17238 (.I0(n7022), .I1(n2630), .I2(n11232), .O(n7051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17238.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17239 (.I0(n2597), .I1(n6989), .I2(n11181), .O(n7020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17239.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17240 (.I0(n7020), .I1(n2628), .I2(n11232), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17240.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17241 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n7051), 
            .I2(n11254), .O(n11255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__17241.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__17242 (.I0(n2601), .I1(n6993), .I2(n11181), .O(n7024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17242.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17243 (.I0(n7024), .I1(n2632), .I2(n11232), .O(n7053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17243.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17244 (.I0(n2603), .I1(n6995), .I2(n11181), .O(n7026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17244.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17245 (.I0(n7026), .I1(n2634), .I2(n11232), .O(n7055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17245.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17246 (.I0(n7055), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n7053), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17246.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17247 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7057), 
            .I2(n11255), .I3(n11256), .O(n11257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__17247.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__17248 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n7053), .I3(n7055), .O(n11258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17248.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17249 (.I0(n7051), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n11254), .O(n11259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17249.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17250 (.I0(n7020), .I1(n2628), .I2(n11232), .O(n7049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17250.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17251 (.I0(n7049), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n7051), 
            .O(n11260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17251.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17252 (.I0(n2595), .I1(n6987), .I2(n11181), .O(n7018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17252.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17253 (.I0(n7018), .I1(n2626), .I2(n11232), .O(n7047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17253.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17254 (.I0(n7016), .I1(n2624), .I2(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I3(n11232), .O(n11261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17254.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17255 (.I0(n2592), .I1(n6983), .I2(n11181), .O(n7014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17255.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17256 (.I0(n7014), .I1(n2623), .I2(n11232), .I3(n9976), 
            .O(n11262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__17256.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__17257 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n7047), 
            .I2(n11261), .I3(n11262), .O(n11263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__17257.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__17258 (.I0(n11259), .I1(n11258), .I2(n11260), .I3(n11263), 
            .O(n11264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__17258.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__17259 (.I0(n11248), .I1(n11253), .I2(n11257), .I3(n11264), 
            .O(n11265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17259.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17260 (.I0(n7833), .I1(n7047), .I2(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[15] ), .O(n11266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17260.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17261 (.I0(n7014), .I1(n2623), .I2(n11232), .O(n7831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17261.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17262 (.I0(n11266), .I1(n7831), .I2(n9976), .O(n11267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8e8 */ ;
    defparam LUT__17262.LUTMASK = 16'he8e8;
    EFX_LUT4 LUT__17263 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n11267), 
            .I2(n10091), .O(n11268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17263.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17264 (.I0(n11265), .I1(n11268), .O(n11269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17264.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17265 (.I0(n7833), .I1(n3414), .I2(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I3(n11269), .O(n11270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17265.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17266 (.I0(n7831), .I1(n3413), .I2(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I3(n11269), .O(n11271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17266.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17267 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n7831), 
            .I2(n10091), .O(n11272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17267.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17268 (.I0(n11271), .I1(n11270), .I2(n11272), .O(n11273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__17268.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__17269 (.I0(n3414), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n2656), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17269.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17270 (.I0(n7833), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n7047), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17270.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17271 (.I0(n11275), .I1(n11274), .I2(n11269), .I3(n11272), 
            .O(n11276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__17271.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__17272 (.I0(n11273), .I1(n11276), .I2(\u_black_pixel_avg/y_sum[13] ), 
            .O(n11277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17272.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17273 (.I0(n2686), .I1(\u_black_pixel_avg/y_sum[14] ), 
            .I2(n11265), .I3(n11268), .O(n7104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17273.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17274 (.I0(n7104), .I1(\u_black_pixel_avg/y_sum[13] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17274.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17275 (.I0(\u_black_pixel_avg/y_sum[15] ), .I1(n2654), 
            .I2(n11232), .O(n7075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17275.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17276 (.I0(n7075), .I1(n2684), .I2(n11269), .O(n7102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17276.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17277 (.I0(n7044), .I1(n2652), .I2(n11232), .O(n7073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17277.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17278 (.I0(n2682), .I1(n7073), .I2(n11265), .I3(n11268), 
            .O(n7100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17278.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17279 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n2678), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n2680), .O(n11279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17279.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17280 (.I0(n2676), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n11279), .O(n11280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17280.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17281 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n7069), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n7071), .O(n11281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17281.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17282 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n7067), 
            .I2(n11281), .O(n11282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17282.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17283 (.I0(n11280), .I1(n11282), .I2(n11265), .I3(n11268), 
            .O(n11283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17283.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17284 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n7100), 
            .I2(n11283), .O(n11284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17284.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17285 (.I0(n11278), .I1(n7102), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n11284), .O(n11285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__17285.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__17286 (.I0(n2678), .I1(n7069), .I2(n11265), .I3(n11268), 
            .O(n7096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17286.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17287 (.I0(n2676), .I1(n7067), .I2(n11265), .I3(n11268), 
            .O(n7094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17287.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17288 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n7094), 
            .I2(n7096), .I3(\u_black_pixel_avg/black_pixel_count[5] ), .O(n11286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17288.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17289 (.I0(n2680), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n2682), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n11287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17289.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17290 (.I0(n7073), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n7071), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17290.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17291 (.I0(n11288), .I1(n11287), .I2(n11269), .I3(n11283), 
            .O(n11289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17291.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17292 (.I0(n7065), .I1(n2674), .I2(n11269), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17292.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17293 (.I0(n11289), .I1(n11290), .I2(n11286), .O(n11291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17293.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17294 (.I0(n2668), .I1(n7059), .I2(n11265), .I3(n11268), 
            .O(n7086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17294.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17295 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7086), 
            .O(n11292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17295.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17296 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n2664), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n2666), 
            .O(n11293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17296.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17297 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n2656), 
            .O(n11294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17297.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17298 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n2658), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n2660), 
            .O(n11295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17298.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17299 (.I0(n2662), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n11294), .I3(n11295), .O(n11296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17299.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17300 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n7049), 
            .O(n11297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17300.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17301 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n7047), 
            .O(n11298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17301.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17302 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n7053), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n7051), 
            .O(n11299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17302.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17303 (.I0(n11297), .I1(n11298), .I2(n11299), .O(n11300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17303.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17304 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7055), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n7057), 
            .O(n11301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17304.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17305 (.I0(n11300), .I1(n11301), .O(n11302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17305.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17306 (.I0(n11296), .I1(n11293), .I2(n11302), .I3(n11269), 
            .O(n11303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__17306.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__17307 (.I0(n7065), .I1(n2674), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11269), .O(n11304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17307.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17308 (.I0(n2670), .I1(n7061), .I2(n11265), .I3(n11268), 
            .O(n7088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17308.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17309 (.I0(n7034), .I1(n2642), .I2(n11232), .O(n7063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17309.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17310 (.I0(n2672), .I1(n7063), .I2(n11265), .I3(n11268), 
            .O(n7090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17310.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17311 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n7090), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7088), .O(n11305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17311.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17312 (.I0(n11292), .I1(n11303), .I2(n11304), .I3(n11305), 
            .O(n11306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__17312.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__17313 (.I0(n11291), .I1(n11285), .I2(n11273), .I3(n11306), 
            .O(n11307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17313.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17314 (.I0(n7088), .I1(n7090), .I2(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17314.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17315 (.I0(n2666), .I1(n7057), .I2(n11265), .I3(n11268), 
            .O(n7084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17315.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17316 (.I0(n7084), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n7086), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17316.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17317 (.I0(n11292), .I1(n11308), .I2(n11309), .I3(n11303), 
            .O(n11310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__17317.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__17318 (.I0(n2660), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n2658), .O(n11311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17318.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17319 (.I0(n11311), .I1(n7049), .I2(n11268), .O(n11312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__17319.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__17320 (.I0(n2658), .I1(n2660), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17320.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17321 (.I0(n11297), .I1(n7051), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17321.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17322 (.I0(n11313), .I1(n11314), .I2(n11265), .I3(n11268), 
            .O(n11315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17322.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17323 (.I0(n11294), .I1(n11298), .I2(n11265), .I3(n11268), 
            .O(n11316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17323.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17324 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n11312), 
            .I2(n11315), .I3(n11316), .O(n11317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__17324.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__17325 (.I0(n2662), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n2664), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17325.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17326 (.I0(n7055), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n7053), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n11319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17326.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17327 (.I0(n11319), .I1(n11300), .O(n11320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17327.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17328 (.I0(n11318), .I1(n11296), .I2(n11320), .I3(n11269), 
            .O(n11321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__17328.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__17329 (.I0(n11317), .I1(n11276), .I2(n11321), .O(n11322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17329.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17330 (.I0(n11322), .I1(n11310), .I2(n11273), .O(n11323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__17330.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__17331 (.I0(n11307), .I1(n11323), .O(n11324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__17331.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__17332 (.I0(n11270), .I1(n11271), .I2(\u_black_pixel_avg/y_sum[13] ), 
            .O(n11325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17332.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17333 (.I0(n11310), .I1(n11317), .I2(n11321), .I3(n11325), 
            .O(n11326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__17333.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__17334 (.I0(n11291), .I1(n11285), .I2(n11306), .I3(n11325), 
            .O(n11327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__17334.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__17335 (.I0(n2716), .I1(n11324), .I2(n11326), .I3(n11327), 
            .O(n11328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__17335.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__17336 (.I0(n11277), .I1(n11328), .O(n7131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__17336.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__17337 (.I0(\u_black_pixel_avg/y_sum[12] ), .I1(n9702), 
            .O(n11329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17337.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17338 (.I0(\u_black_pixel_avg/y_sum[12] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17338.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17339 (.I0(n11277), .I1(n11327), .I2(n11326), .I3(n11330), 
            .O(n11331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17339.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17340 (.I0(n2716), .I1(n11324), .I2(n11331), .O(n11332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__17340.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__17341 (.I0(n7104), .I1(n2714), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n11324), .O(n11333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17341.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17342 (.I0(n2712), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n2714), .I3(\u_black_pixel_avg/black_pixel_count[2] ), .O(n11334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17342.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17343 (.I0(n7104), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n7102), .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n11335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17343.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17344 (.I0(n2708), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n2710), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17344.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17345 (.I0(n7071), .I1(n2680), .I2(n11269), .O(n7098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17345.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17346 (.I0(n7100), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n7098), .I3(\u_black_pixel_avg/black_pixel_count[5] ), .O(n11337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17346.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17347 (.I0(n11336), .I1(n11337), .I2(n11307), .I3(n11323), 
            .O(n11338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17347.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17348 (.I0(n11335), .I1(n11334), .I2(n11338), .I3(n11324), 
            .O(n11339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17348.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17349 (.I0(n11332), .I1(n11329), .I2(n11333), .I3(n11339), 
            .O(n11340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__17349.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__17350 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n2710), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n2712), .O(n11341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17350.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17351 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7100), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n7102), .O(n11342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17351.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17352 (.I0(n11342), .I1(n11341), .I2(n11338), .I3(n11324), 
            .O(n11343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17352.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17353 (.I0(n7098), .I1(n2708), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n11324), .O(n11344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17353.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17354 (.I0(n7096), .I1(n2706), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n11324), .O(n11345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17354.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17355 (.I0(n11343), .I1(n11344), .I2(n11345), .O(n11346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__17355.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__17356 (.I0(n7096), .I1(n2706), .I2(n11324), .O(n7121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17356.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17357 (.I0(n2704), .I1(n7094), .I2(n11307), .I3(n11323), 
            .O(n7119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17357.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17358 (.I0(n7119), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17358.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17359 (.I0(n2700), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n2702), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17359.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17360 (.I0(n7065), .I1(n2674), .I2(n11269), .O(n7092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17360.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17361 (.I0(n7090), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n7092), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17361.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17362 (.I0(n2696), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n2698), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17362.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17363 (.I0(n7088), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n7086), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17363.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17364 (.I0(n11350), .I1(n11351), .I2(n11307), .I3(n11323), 
            .O(n11352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17364.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17365 (.I0(n11349), .I1(n11348), .I2(n11352), .I3(n11324), 
            .O(n11353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17365.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17366 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n7121), 
            .I2(n11347), .I3(n11353), .O(n11354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17366.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17367 (.I0(n2702), .I1(n7092), .I2(n11307), .I3(n11323), 
            .O(n7117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__17367.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__17368 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n7117), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n7119), .O(n11355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17368.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17369 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n2690), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n2692), 
            .O(n11356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17369.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17370 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n2694), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n2696), 
            .O(n11357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17370.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17371 (.I0(n7055), .I1(n2664), .I2(n11269), .O(n7082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17371.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17372 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n7086), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n7082), 
            .O(n11358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17372.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17373 (.I0(n7053), .I1(n2662), .I2(n11269), .O(n7080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17373.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17374 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7084), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n7080), 
            .O(n11359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17374.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17375 (.I0(n11358), .I1(n11359), .O(n11360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17375.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17376 (.I0(n11357), .I1(n11356), .I2(n11360), .I3(n11324), 
            .O(n11361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__17376.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__17377 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n2698), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n2700), .O(n11362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17377.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17378 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n7090), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n7088), 
            .O(n11363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17378.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17379 (.I0(n11363), .I1(n11362), .I2(n11352), .I3(n11324), 
            .O(n11364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17379.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17380 (.I0(n11355), .I1(n11353), .I2(n11361), .I3(n11364), 
            .O(n11365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__17380.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__17381 (.I0(n11340), .I1(n11346), .I2(n11354), .I3(n11365), 
            .O(n11366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17381.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17382 (.I0(n7080), .I1(n2690), .I2(n11324), .O(n7821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17382.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17383 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n7821), 
            .O(n11367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17383.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17384 (.I0(n7082), .I1(n2692), .I2(n11324), .O(n7107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17384.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17385 (.I0(n7084), .I1(n2694), .I2(n11324), .O(n7109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17385.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17386 (.I0(n7107), .I1(n7109), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[12] ), .O(n11368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17386.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17387 (.I0(n7051), .I1(n2660), .I2(n11269), .O(n7078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17387.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17388 (.I0(n7078), .I1(n2688), .I2(n11324), .O(n7819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17388.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17389 (.I0(n7819), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n7821), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17389.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17390 (.I0(n7047), .I1(n2656), .I2(n11269), .O(n7827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17390.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17391 (.I0(n7827), .I1(n3409), .I2(n11324), .O(n7815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17391.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17392 (.I0(n7049), .I1(n2658), .I2(n11269), .O(n7829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17392.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17393 (.I0(n7829), .I1(n3411), .I2(n11324), .O(n7817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17393.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17394 (.I0(n7817), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I2(n7815), .I3(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n11370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17394.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17395 (.I0(n11368), .I1(n11367), .I2(n11369), .I3(n11370), 
            .O(n11371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__17395.LUTMASK = 16'he000;
    EFX_LUT4 LUT__17396 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n7817), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n7819), 
            .O(n11372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17396.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17397 (.I0(n7831), .I1(n3413), .I2(n11269), .O(n7823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17397.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17398 (.I0(n7823), .I1(n3406), .I2(n11324), .O(n7811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17398.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17399 (.I0(n7811), .I1(n10091), .O(n11373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17399.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17400 (.I0(n7833), .I1(n3414), .I2(n11269), .O(n7825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17400.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17401 (.I0(n7825), .I1(n3407), .I2(n11324), .O(n7813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17401.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17402 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n7815), 
            .I2(\u_black_pixel_avg/black_pixel_count[18] ), .I3(n7813), 
            .O(n11374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17402.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17403 (.I0(n11372), .I1(n11370), .I2(n11373), .I3(n11374), 
            .O(n11375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__17403.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__17404 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n7823), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(n10090), 
            .O(n11376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17404.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17405 (.I0(n7813), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n11376), .I3(n11373), .O(n11377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__17405.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__17406 (.I0(n11366), .I1(n11371), .I2(n11375), .I3(n11377), 
            .O(n11378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__17406.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__17407 (.I0(n7131), .I1(n2742), .I2(n11378), .O(n7154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17407.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17408 (.I0(\u_black_pixel_avg/y_sum[11] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17408.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17409 (.I0(\u_black_pixel_avg/y_sum[11] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17409.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17410 (.I0(\u_black_pixel_avg/y_sum[12] ), .I1(n2744), 
            .I2(n11380), .I3(n11378), .O(n11381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17410.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17411 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n7154), 
            .I2(n11379), .I3(n11381), .O(n11382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hddd4 */ ;
    defparam LUT__17411.LUTMASK = 16'hddd4;
    EFX_LUT4 LUT__17412 (.I0(n7104), .I1(n2714), .I2(n11324), .O(n7129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17412.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17413 (.I0(n7129), .I1(n2740), .I2(n11378), .O(n7152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17413.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17414 (.I0(n7102), .I1(n2712), .I2(n11324), .O(n7127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17414.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17415 (.I0(n7127), .I1(n2738), .I2(n11378), .O(n7150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17415.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17416 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7150), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n7152), .O(n11383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17416.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17417 (.I0(n7152), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n11382), .I3(n11383), .O(n11384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17417.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17418 (.I0(n7100), .I1(n2710), .I2(n11324), .O(n7125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17418.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17419 (.I0(n7125), .I1(n2736), .I2(n11378), .O(n7148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17419.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17420 (.I0(n7148), .I1(n7150), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17420.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17421 (.I0(n7098), .I1(n2708), .I2(n11324), .O(n7123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17421.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17422 (.I0(n7123), .I1(n2734), .I2(n11378), .O(n7146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17422.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17423 (.I0(n7121), .I1(n2732), .I2(n11378), .O(n7144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17423.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17424 (.I0(n7144), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17424.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17425 (.I0(n11385), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n7146), .I3(n11386), .O(n11387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17425.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17426 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n7146), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n7148), .O(n11388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17426.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17427 (.I0(n7109), .I1(n2720), .I2(n11378), .O(n7764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17427.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17428 (.I0(n7107), .I1(n2718), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I3(n11378), .O(n11389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17428.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17429 (.I0(n7821), .I1(n3404), .I2(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I3(n11378), .O(n11390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17429.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17430 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n7764), 
            .I2(n11389), .I3(n11390), .O(n11391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__17430.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__17431 (.I0(n7086), .I1(n2696), .I2(n11324), .O(n7111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17431.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17432 (.I0(n7111), .I1(n2722), .I2(n11378), .O(n7134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17432.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17433 (.I0(n7088), .I1(n2698), .I2(n11324), .O(n7113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17433.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17434 (.I0(n7113), .I1(n2724), .I2(n11378), .O(n7136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17434.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17435 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n7136), 
            .I2(\u_black_pixel_avg/black_pixel_count[12] ), .I3(n7134), 
            .O(n11392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17435.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17436 (.I0(n7119), .I1(n2730), .I2(n11378), .O(n7142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17436.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17437 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n7142), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n7144), .O(n11393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17437.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17438 (.I0(n7117), .I1(n2728), .I2(n11378), .O(n7140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17438.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17439 (.I0(n7090), .I1(n2700), .I2(n11324), .O(n7115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17439.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17440 (.I0(n7115), .I1(n2726), .I2(n11378), .O(n7138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17440.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17441 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7138), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7140), .O(n11394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17441.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17442 (.I0(n11391), .I1(n11392), .I2(n11393), .I3(n11394), 
            .O(n11395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__17442.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__17443 (.I0(n11384), .I1(n11388), .I2(n11387), .I3(n11395), 
            .O(n11396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__17443.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__17444 (.I0(n11391), .I1(n11392), .O(n11397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17444.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17445 (.I0(n7140), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n7142), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17445.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17446 (.I0(n7138), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n7136), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17446.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17447 (.I0(n11398), .I1(n11394), .I2(n11399), .O(n11400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17447.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17448 (.I0(n7134), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n7764), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n11401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17448.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17449 (.I0(n11401), .I1(n11391), .O(n11402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17449.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17450 (.I0(n7107), .I1(n2718), .I2(n11378), .O(n7762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17450.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17451 (.I0(n7762), .I1(n11390), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17451.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17452 (.I0(n7821), .I1(n3404), .I2(n11378), .O(n7760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17452.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17453 (.I0(n7817), .I1(n3400), .I2(n11378), .O(n7756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17453.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17454 (.I0(n7756), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n7760), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n11404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17454.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17455 (.I0(n7819), .I1(n3402), .I2(n11378), .O(n7758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17455.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17456 (.I0(n7815), .I1(n3398), .I2(n11378), .O(n7754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17456.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17457 (.I0(n7754), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n7758), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17457.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17458 (.I0(n11403), .I1(n11404), .I2(n11405), .O(n11406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17458.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17459 (.I0(n11400), .I1(n11397), .I2(n11402), .I3(n11406), 
            .O(n11407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__17459.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__17460 (.I0(n7813), .I1(n3396), .I2(n11378), .O(n7752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17460.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17461 (.I0(n7811), .I1(n3395), .I2(n11378), .O(n7750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17461.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17462 (.I0(\u_black_pixel_avg/black_pixel_count[20] ), .I1(n7750), 
            .O(n11408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17462.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17463 (.I0(n7756), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[16] ), .I3(n7758), 
            .O(n11409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17463.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17464 (.I0(n11409), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n7754), .O(n11410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__17464.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__17465 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n7752), 
            .I2(n11408), .I3(n11410), .O(n11411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__17465.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__17466 (.I0(n7750), .I1(n7752), .I2(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[19] ), .O(n11412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17466.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17467 (.I0(n11412), .I1(n10090), .O(n11413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17467.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17468 (.I0(n11396), .I1(n11407), .I2(n11411), .I3(n11413), 
            .O(n11414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17468.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17469 (.I0(n7154), .I1(n2766), .I2(n11414), .O(n7201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17469.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17470 (.I0(\u_black_pixel_avg/y_sum[11] ), .I1(n2770), 
            .I2(n11414), .O(n7205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17470.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17471 (.I0(n7205), .I1(\u_black_pixel_avg/y_sum[10] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17471.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17472 (.I0(\u_black_pixel_avg/y_sum[12] ), .I1(n2744), 
            .I2(n11378), .O(n7156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17472.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17473 (.I0(n7156), .I1(n2768), .I2(n11414), .O(n7203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17473.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17474 (.I0(n7152), .I1(n2764), .I2(n11414), .O(n7199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17474.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17475 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n7201), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n7199), .O(n11416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17475.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17476 (.I0(n11415), .I1(n7203), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I3(n11416), .O(n11417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__17476.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__17477 (.I0(n7144), .I1(n2756), .I2(n11414), .O(n7191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17477.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17478 (.I0(n7142), .I1(n2754), .I2(n11414), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17478.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17479 (.I0(n7146), .I1(n2758), .I2(n11414), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17479.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17480 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n7191), 
            .I2(n11418), .I3(n11419), .O(n11420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__17480.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__17481 (.I0(n7148), .I1(n2760), .I2(n11414), .O(n7195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17481.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17482 (.I0(n7150), .I1(n2762), .I2(n11414), .O(n7197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17482.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17483 (.I0(n7197), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n7195), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n11421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17483.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17484 (.I0(n7199), .I1(n7201), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n11422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17484.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17485 (.I0(n11420), .I1(n11421), .I2(n11422), .O(n11423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__17485.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__17486 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n7197), 
            .O(n11424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17486.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17487 (.I0(n11424), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I2(n7195), .I3(n11420), .O(n11425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__17487.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__17488 (.I0(n7146), .I1(n2758), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11414), .O(n11426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17488.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17489 (.I0(n7191), .I1(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I2(n11426), .I3(n11418), .O(n11427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17489.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17490 (.I0(n7138), .I1(n2750), .I2(n11414), .O(n7185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17490.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17491 (.I0(n7136), .I1(n2748), .I2(n11414), .O(n7748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17491.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17492 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7748), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n7185), 
            .O(n11428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17492.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17493 (.I0(n7134), .I1(n2746), .I2(n11414), .O(n7746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17493.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17494 (.I0(n7764), .I1(n3348), .I2(n11414), .O(n7744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17494.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17495 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n7744), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n7746), 
            .O(n11429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17495.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17496 (.I0(n7142), .I1(n2754), .I2(n11414), .O(n7189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17496.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17497 (.I0(n7140), .I1(n2752), .I2(n11414), .O(n7187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17497.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17498 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7187), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7189), .O(n11430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17498.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17499 (.I0(n11427), .I1(n11428), .I2(n11429), .I3(n11430), 
            .O(n11431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__17499.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__17500 (.I0(n11423), .I1(n11417), .I2(n11425), .I3(n11431), 
            .O(n11432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17500.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17501 (.I0(n7187), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n7185), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17501.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17502 (.I0(n7746), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n7748), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17502.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17503 (.I0(n11433), .I1(n11428), .I2(n11434), .I3(n11429), 
            .O(n11435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17503.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17504 (.I0(n7754), .I1(n3338), .I2(n11414), .O(n7729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17504.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17505 (.I0(n7756), .I1(n3340), .I2(n11414), .O(n7731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17505.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17506 (.I0(n7731), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n7729), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n11436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17506.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17507 (.I0(n7760), .I1(n3344), .I2(n11414), .O(n7735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17507.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17508 (.I0(n7758), .I1(n3342), .I2(n11414), .O(n7733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17508.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17509 (.I0(n7733), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n7735), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17509.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17510 (.I0(n11436), .I1(n11437), .O(n11438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17510.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17511 (.I0(n7762), .I1(n3346), .I2(n11414), .O(n7742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17511.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17512 (.I0(n7744), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n7742), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n11439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17512.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17513 (.I0(n11435), .I1(n11438), .I2(n11439), .O(n11440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17513.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17514 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n7742), 
            .I2(\u_black_pixel_avg/black_pixel_count[16] ), .I3(n7735), 
            .O(n11441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17514.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17515 (.I0(n7731), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n7733), 
            .O(n11442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17515.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17516 (.I0(n11442), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I2(n7729), .O(n11443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__17516.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__17517 (.I0(n7750), .I1(n3335), .I2(n11414), .O(n7725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17517.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17518 (.I0(n7752), .I1(n3336), .I2(n11414), .O(n7727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17518.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17519 (.I0(\u_black_pixel_avg/black_pixel_count[20] ), .I1(n7727), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(n7725), 
            .O(n11444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17519.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17520 (.I0(n11441), .I1(n11438), .I2(n11443), .I3(n11444), 
            .O(n11445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__17520.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__17521 (.I0(n7725), .I1(n7727), .I2(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[20] ), .O(n11446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17521.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17522 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n10251), 
            .I2(n11446), .O(n11447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17522.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17523 (.I0(n11432), .I1(n11440), .I2(n11445), .I3(n11447), 
            .O(n11448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17523.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17524 (.I0(n7201), .I1(n2804), .I2(n11448), .O(n7257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17524.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17525 (.I0(n7203), .I1(n2806), .I2(n11448), .O(n7259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17525.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17526 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n7259), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n7257), .O(n11449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17526.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17527 (.I0(n7205), .I1(n2808), .I2(n11448), .O(n7261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17527.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17528 (.I0(\u_black_pixel_avg/y_sum[9] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17528.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17529 (.I0(\u_black_pixel_avg/y_sum[9] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17529.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17530 (.I0(\u_black_pixel_avg/y_sum[10] ), .I1(n2810), 
            .I2(n11451), .I3(n11448), .O(n11452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17530.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17531 (.I0(n7261), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n11450), .I3(n11452), .O(n11453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hddd4 */ ;
    defparam LUT__17531.LUTMASK = 16'hddd4;
    EFX_LUT4 LUT__17532 (.I0(n7199), .I1(n2802), .I2(n11448), .O(n7255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17532.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17533 (.I0(n7255), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n11454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17533.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17534 (.I0(n7257), .I1(n7259), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[3] ), .O(n11455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17534.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17535 (.I0(n11453), .I1(n11449), .I2(n11454), .I3(n11455), 
            .O(n11456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__17535.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__17536 (.I0(n7748), .I1(n3333), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n11448), .O(n11457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17536.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17537 (.I0(n7746), .I1(n3331), .I2(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I3(n11448), .O(n11458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17537.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17538 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n3317), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n3319), 
            .O(n11459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17538.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17539 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n7733), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n7735), 
            .O(n11460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17539.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17540 (.I0(n11460), .I1(n11459), .I2(n11448), .O(n11461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17540.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17541 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n3327), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n3329), 
            .O(n11462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17541.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17542 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n7744), 
            .I2(\u_black_pixel_avg/black_pixel_count[16] ), .I3(n7742), 
            .O(n11463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17542.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17543 (.I0(n11463), .I1(n11462), .I2(n11448), .O(n11464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17543.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17544 (.I0(n11457), .I1(n11458), .I2(n11461), .I3(n11464), 
            .O(n11465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17544.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17545 (.I0(n7187), .I1(n2790), .I2(n11448), .O(n7723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17545.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17546 (.I0(n7185), .I1(n2788), .I2(n11448), .O(n7721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17546.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17547 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7721), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n7723), 
            .O(n11466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17547.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17548 (.I0(n7191), .I1(n2794), .I2(n11448), .O(n7247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17548.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17549 (.I0(n7189), .I1(n2792), .I2(n11448), .O(n7245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17549.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17550 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7245), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7247), .O(n11467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17550.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17551 (.I0(n11465), .I1(n11466), .I2(n11467), .O(n11468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__17551.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__17552 (.I0(n7195), .I1(n2798), .I2(n11448), .O(n7251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17552.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17553 (.I0(n7146), .I1(n2758), .I2(n11414), .O(n7193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17553.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17554 (.I0(n7193), .I1(n2796), .I2(n11448), .O(n7249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17554.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17555 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n7249), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n7251), .O(n11469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17555.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17556 (.I0(n7197), .I1(n2800), .I2(n11448), .O(n7253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17556.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17557 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n7253), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n7255), .O(n11470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17557.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17558 (.I0(n11456), .I1(n11468), .I2(n11469), .I3(n11470), 
            .O(n11471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__17558.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__17559 (.I0(n7251), .I1(n7253), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n11472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17559.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17560 (.I0(n11472), .I1(n7249), .I2(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n11473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__17560.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__17561 (.I0(n7247), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n11473), .I3(n11468), .O(n11474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__17561.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__17562 (.I0(n7746), .I1(n3331), .I2(n11448), .O(n7717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17562.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17563 (.I0(n7744), .I1(n3329), .I2(n11448), .O(n7715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17563.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17564 (.I0(n7715), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n7717), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17564.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17565 (.I0(n7735), .I1(n3319), .I2(n11448), .O(n7711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17565.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17566 (.I0(n7742), .I1(n3327), .I2(n11448), .O(n7713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17566.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17567 (.I0(n7713), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I2(n7711), .I3(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n11476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17567.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17568 (.I0(n11464), .I1(n11475), .I2(n11476), .I3(n11461), 
            .O(n11477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__17568.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__17569 (.I0(n7245), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(n7723), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17569.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17570 (.I0(n7748), .I1(n3333), .I2(n11448), .O(n7719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17570.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17571 (.I0(n7721), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I2(n7719), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n11479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17571.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17572 (.I0(n11478), .I1(n11466), .I2(n11479), .I3(n11465), 
            .O(n11480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17572.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17573 (.I0(n7729), .I1(n3313), .I2(n11448), .O(n7705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17573.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17574 (.I0(n7727), .I1(n3311), .I2(n11448), .O(n7703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17574.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17575 (.I0(n7703), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I2(n7705), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n11481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17575.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17576 (.I0(n7725), .I1(n3310), .I2(n11448), .O(n7701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17576.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17577 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n7701), 
            .I2(n10251), .O(n11482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17577.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17578 (.I0(n7731), .I1(n3315), .I2(n11448), .O(n7707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17578.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17579 (.I0(n7733), .I1(n3317), .I2(n11448), .O(n7709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17579.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17580 (.I0(n7709), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n7707), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n11483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17580.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17581 (.I0(n11481), .I1(n11482), .I2(n11483), .O(n11484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__17581.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__17582 (.I0(n11477), .I1(n11480), .I2(n11484), .O(n11485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__17582.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__17583 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n7707), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(n7705), 
            .O(n11486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17583.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17584 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n7701), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(n7703), 
            .O(n11487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17584.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17585 (.I0(n11486), .I1(n11481), .I2(n11487), .I3(n11482), 
            .O(n11488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17585.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17586 (.I0(n11474), .I1(n11471), .I2(n11485), .I3(n11488), 
            .O(n11489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__17586.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__17587 (.I0(n10853), .I1(n10852), .I2(n11489), .O(n11490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17587.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17588 (.I0(\u_black_pixel_avg/y_sum[10] ), .I1(n2810), 
            .I2(n11448), .O(n7263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17588.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17589 (.I0(n2860), .I1(n7263), .I2(n11489), .O(n7348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17589.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17590 (.I0(n2858), .I1(n7261), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n11491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17590.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17591 (.I0(n11490), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n7348), .I3(n11491), .O(n11492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17591.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17592 (.I0(n2858), .I1(n7261), .I2(n11489), .O(n7346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17592.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17593 (.I0(n2856), .I1(n7259), .I2(n11489), .O(n7344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17593.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17594 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7344), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n7346), .O(n11493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17594.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17595 (.I0(n2854), .I1(n7257), .I2(n11489), .O(n7342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17595.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17596 (.I0(n7342), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n7344), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17596.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17597 (.I0(n2848), .I1(n7251), .I2(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I3(n11489), .O(n11495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17597.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17598 (.I0(n2850), .I1(n7253), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11489), .O(n11496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17598.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17599 (.I0(n2854), .I1(n7257), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n11489), .O(n11497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17599.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17600 (.I0(n2852), .I1(n7255), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n11489), .O(n11498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17600.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17601 (.I0(n11495), .I1(n11496), .I2(n11497), .I3(n11498), 
            .O(n11499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17601.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17602 (.I0(n11492), .I1(n11493), .I2(n11494), .I3(n11499), 
            .O(n11500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17602.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17603 (.I0(n2850), .I1(n7253), .I2(n11489), .O(n7338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17603.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17604 (.I0(n2852), .I1(n7255), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17604.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17605 (.I0(n7338), .I1(n11501), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11495), .O(n11502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__17605.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__17606 (.I0(n2848), .I1(n7251), .I2(n11489), .O(n7336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17606.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17607 (.I0(n2846), .I1(n7249), .I2(n11489), .O(n7334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17607.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17608 (.I0(n7334), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n7336), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17608.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17609 (.I0(n2844), .I1(n7247), .I2(n11489), .O(n7692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17609.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17610 (.I0(n2842), .I1(n7245), .I2(n11489), .O(n7690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17610.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17611 (.I0(n7690), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n7692), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17611.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17612 (.I0(n11502), .I1(n11503), .I2(n11504), .O(n11505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17612.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17613 (.I0(n7692), .I1(\u_black_pixel_avg/black_pixel_count[10] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7334), .O(n11506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17613.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17614 (.I0(n3308), .I1(n7723), .I2(n11489), .O(n7688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17614.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17615 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7688), 
            .O(n11507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17615.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17616 (.I0(n11506), .I1(n7690), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(n11507), .O(n11508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17616.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17617 (.I0(n3298), .I1(n7713), .I2(n11489), .O(n7678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17617.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17618 (.I0(n3300), .I1(n7715), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17618.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17619 (.I0(n3296), .I1(n7711), .I2(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I3(n11489), .O(n11510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17619.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17620 (.I0(n7678), .I1(n11509), .I2(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I3(n11510), .O(n11511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__17620.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__17621 (.I0(n3290), .I1(n7705), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[21] ), 
            .O(n11512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17621.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17622 (.I0(n3292), .I1(n7707), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n11513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17622.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17623 (.I0(n3294), .I1(n7709), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n11514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17623.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17624 (.I0(n3296), .I1(n7711), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n11515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17624.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17625 (.I0(n11512), .I1(n11513), .I2(n11514), .I3(n11515), 
            .O(n11516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17625.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17626 (.I0(n3302), .I1(n7717), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n11517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17626.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17627 (.I0(n3304), .I1(n7719), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17627.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17628 (.I0(n3306), .I1(n7721), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n11519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17628.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17629 (.I0(n3308), .I1(n7723), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17629.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17630 (.I0(n11517), .I1(n11518), .I2(n11519), .I3(n11520), 
            .O(n11521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17630.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17631 (.I0(n3288), .I1(n7703), .I2(n11489), .O(n7668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17631.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17632 (.I0(n3287), .I1(n7701), .I2(n11489), .I3(\u_black_pixel_avg/black_pixel_count[23] ), 
            .O(n11522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17632.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17633 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n7668), 
            .I2(n11522), .I3(n10250), .O(n11523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17633.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17634 (.I0(n11511), .I1(n11516), .I2(n11521), .I3(n11523), 
            .O(n11524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__17634.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__17635 (.I0(n11500), .I1(n11505), .I2(n11508), .I3(n11524), 
            .O(n11525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17635.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17636 (.I0(n3304), .I1(n7719), .I2(n11489), .O(n7684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17636.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17637 (.I0(n3306), .I1(n7721), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n11489), .O(n11526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17637.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17638 (.I0(n7684), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n11526), .I3(n11517), .O(n11527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17638.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17639 (.I0(n3298), .I1(n7713), .I2(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I3(n11489), .O(n11528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17639.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17640 (.I0(n3302), .I1(n7717), .I2(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I3(n11489), .O(n11529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17640.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17641 (.I0(n3300), .I1(n7715), .I2(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I3(n11489), .O(n11530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17641.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17642 (.I0(n11510), .I1(n11528), .I2(n11529), .I3(n11530), 
            .O(n11531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17642.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17643 (.I0(n11531), .I1(n11527), .I2(n11511), .I3(n11516), 
            .O(n11532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17643.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17644 (.I0(n3292), .I1(n7707), .I2(n11489), .O(n7672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17644.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17645 (.I0(n3294), .I1(n7709), .I2(n11489), .O(n7674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17645.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17646 (.I0(n7672), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[19] ), .I3(n7674), 
            .O(n11533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17646.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17647 (.I0(n3290), .I1(n7705), .I2(n11489), .O(n7670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17647.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17648 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n7668), 
            .O(n11534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17648.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17649 (.I0(n11533), .I1(n7670), .I2(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I3(n11534), .O(n11535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17649.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17650 (.I0(n3287), .I1(n7701), .I2(n11489), .O(n7666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17650.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17651 (.I0(n7666), .I1(n10251), .O(n11536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17651.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17652 (.I0(n11532), .I1(n11535), .I2(n11523), .I3(n11536), 
            .O(n11537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__17652.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__17653 (.I0(n11525), .I1(n11537), .O(n11538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17653.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17654 (.I0(n2937), .I1(\u_black_pixel_avg/y_sum[8] ), 
            .I2(n11538), .O(n7421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17654.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17655 (.I0(n2933), .I1(n7348), .I2(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I3(n11538), .O(n11539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17655.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17656 (.I0(n7346), .I1(n2931), .I2(n11525), .I3(n11537), 
            .O(n7415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17656.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17657 (.I0(n2862), .I1(\u_black_pixel_avg/y_sum[9] ), 
            .I2(n11489), .O(n7350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17657.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17658 (.I0(\u_black_pixel_avg/y_sum[8] ), .I1(\u_black_pixel_avg/y_sum[7] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17658.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17659 (.I0(n7350), .I1(n11540), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n11541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__17659.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__17660 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n7348), 
            .I2(n11541), .O(n11542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__17660.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__17661 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n2937), 
            .I2(\u_black_pixel_avg/y_sum[7] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17661.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17662 (.I0(n2933), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n11544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17662.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17663 (.I0(n11543), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n2935), .I3(n11544), .O(n11545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17663.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17664 (.I0(n11542), .I1(n11545), .I2(n11525), .I3(n11537), 
            .O(n11546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17664.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17665 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7415), 
            .I2(n11546), .O(n11547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17665.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17666 (.I0(n7344), .I1(n2929), .I2(n11525), .I3(n11537), 
            .O(n7413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17666.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17667 (.I0(n7413), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n7415), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17667.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17668 (.I0(n7342), .I1(n2927), .I2(n11525), .I3(n11537), 
            .O(n7411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17668.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17669 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n7411), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n7413), .O(n11549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17669.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17670 (.I0(n11539), .I1(n11547), .I2(n11548), .I3(n11549), 
            .O(n11550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17670.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17671 (.I0(n7411), .I1(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17671.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17672 (.I0(n2852), .I1(n7255), .I2(n11489), .O(n7340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17672.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17673 (.I0(n7340), .I1(n2925), .I2(n11525), .I3(n11537), 
            .O(n7409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17673.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17674 (.I0(n7409), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17674.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17675 (.I0(n7334), .I1(n2919), .I2(n11525), .I3(n11537), 
            .O(n7653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17675.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17676 (.I0(n7692), .I1(n3277), .I2(n11525), .I3(n11537), 
            .O(n7651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17676.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17677 (.I0(n7651), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n7653), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17677.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17678 (.I0(n7338), .I1(n2923), .I2(n11525), .I3(n11537), 
            .O(n7407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17678.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17679 (.I0(n7336), .I1(n2921), .I2(n11525), .I3(n11537), 
            .O(n7655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17679.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17680 (.I0(n7655), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n7407), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17680.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17681 (.I0(n11551), .I1(n11552), .I2(n11553), .I3(n11554), 
            .O(n11555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__17681.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__17682 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n7407), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n7409), .O(n11556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17682.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17683 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n7655), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n7653), 
            .O(n11557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17683.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17684 (.I0(n11556), .I1(n11554), .I2(n11557), .I3(n11553), 
            .O(n11558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17684.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17685 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n7651), 
            .O(n11559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17685.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17686 (.I0(n3275), .I1(n7690), .I2(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I3(n11538), .O(n11560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17686.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17687 (.I0(n7688), .I1(n3273), .I2(n11525), .I3(n11537), 
            .O(n7647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17687.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17688 (.I0(n3306), .I1(n7721), .I2(n11489), .O(n7686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17688.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17689 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n7686), 
            .O(n11561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17689.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17690 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n3271), 
            .O(n11562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17690.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17691 (.I0(n11561), .I1(n11562), .I2(n11525), .I3(n11537), 
            .O(n11563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17691.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17692 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n7647), 
            .I2(n11563), .O(n11564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17692.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17693 (.I0(n7684), .I1(n3269), .I2(n11525), .I3(n11537), 
            .O(n7643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17693.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17694 (.I0(n3302), .I1(n7717), .I2(n11489), .O(n7682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17694.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17695 (.I0(n7682), .I1(n3267), .I2(n11525), .I3(n11537), 
            .O(n7641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17695.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17696 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n7641), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n7643), 
            .O(n11565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17696.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17697 (.I0(n11559), .I1(n11560), .I2(n11564), .I3(n11565), 
            .O(n11566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__17697.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__17698 (.I0(n11555), .I1(n11550), .I2(n11558), .I3(n11566), 
            .O(n11567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17698.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17699 (.I0(n7643), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n11568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17699.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17700 (.I0(n7686), .I1(n3271), .I2(n11525), .I3(n11537), 
            .O(n7645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17700.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17701 (.I0(n7645), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17701.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17702 (.I0(n7690), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17702.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17703 (.I0(n3275), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17703.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17704 (.I0(n11570), .I1(n11571), .I2(n11525), .I3(n11537), 
            .O(n11572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17704.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17705 (.I0(n7647), .I1(n11572), .I2(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I3(n11563), .O(n11573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__17705.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__17706 (.I0(n11569), .I1(n11573), .I2(n11568), .I3(n11565), 
            .O(n11574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__17706.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__17707 (.I0(n3255), .I1(n7670), .I2(n11538), .I3(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n11575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17707.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17708 (.I0(n11535), .I1(n11532), .I2(n11523), .O(n11576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17708.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17709 (.I0(n7668), .I1(n3253), .I2(n11525), .I3(n11576), 
            .O(n11577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__17709.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__17710 (.I0(n11577), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .O(n11578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__17710.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__17711 (.I0(n11532), .I1(n11535), .I2(n11523), .I3(n10251), 
            .O(n11579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__17711.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__17712 (.I0(n11532), .I1(n11535), .I2(n11523), .I3(n7666), 
            .O(n11580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__17712.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__17713 (.I0(n11579), .I1(n3252), .I2(n11525), .I3(n11580), 
            .O(n7625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc0ce */ ;
    defparam LUT__17713.LUTMASK = 16'hc0ce;
    EFX_LUT4 LUT__17714 (.I0(n7668), .I1(n3253), .I2(n11525), .I3(n11537), 
            .O(n7627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17714.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17715 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(n7627), 
            .I2(\u_black_pixel_avg/black_pixel_count[24] ), .I3(n7625), 
            .O(n11581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17715.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17716 (.I0(\u_black_pixel_avg/black_pixel_count[24] ), .I1(n7666), 
            .I2(\u_black_pixel_avg/black_pixel_count[25] ), .I3(n10089), 
            .O(n11582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17716.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17717 (.I0(n11578), .I1(n11575), .I2(n11581), .I3(n11582), 
            .O(n11583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__17717.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__17718 (.I0(n3300), .I1(n7715), .I2(n11489), .O(n7680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17718.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17719 (.I0(n7680), .I1(n3265), .I2(n11525), .I3(n11537), 
            .O(n7639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17719.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17720 (.I0(n7639), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n11584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17720.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17721 (.I0(n7641), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17721.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17722 (.I0(n7674), .I1(n3259), .I2(n11525), .I3(n11537), 
            .O(n7633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17722.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17723 (.I0(n7672), .I1(n3257), .I2(n11525), .I3(n11537), 
            .O(n7631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17723.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17724 (.I0(n7631), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I2(n7633), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n11586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17724.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17725 (.I0(n7678), .I1(n3263), .I2(n11525), .I3(n11537), 
            .O(n7637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17725.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17726 (.I0(n3296), .I1(n7711), .I2(n11489), .O(n7676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17726.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17727 (.I0(n7676), .I1(n3261), .I2(n11525), .I3(n11537), 
            .O(n7635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17727.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17728 (.I0(n7635), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I2(n7637), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n11587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17728.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17729 (.I0(n11584), .I1(n11585), .I2(n11586), .I3(n11587), 
            .O(n11588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__17729.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__17730 (.I0(n11574), .I1(n11583), .I2(n11588), .O(n11589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17730.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17731 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n7639), 
            .I2(\u_black_pixel_avg/black_pixel_count[18] ), .I3(n7637), 
            .O(n11590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17731.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17732 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n7635), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(n7633), 
            .O(n11591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17732.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17733 (.I0(n11590), .I1(n11587), .I2(n11591), .I3(n11586), 
            .O(n11592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17733.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17734 (.I0(n3255), .I1(n7670), .I2(\u_black_pixel_avg/black_pixel_count[22] ), 
            .I3(n11538), .O(n11593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17734.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17735 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n7631), 
            .I2(n11593), .I3(n11581), .O(n11594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__17735.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__17736 (.I0(n11594), .I1(n11592), .I2(n11583), .O(n11595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17736.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17737 (.I0(n11589), .I1(n11567), .I2(n11595), .O(n11596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__17737.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__17738 (.I0(n3006), .I1(n7421), .I2(n11596), .O(n7486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17738.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17739 (.I0(\u_black_pixel_avg/y_sum[6] ), .I1(n9702), 
            .O(n11597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17739.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17740 (.I0(n3008), .I1(\u_black_pixel_avg/y_sum[7] ), 
            .I2(n11597), .I3(n11596), .O(n11598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17740.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17741 (.I0(\u_black_pixel_avg/y_sum[6] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17741.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17742 (.I0(n7486), .I1(n11598), .I2(n11599), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n11600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8fe */ ;
    defparam LUT__17742.LUTMASK = 16'ha8fe;
    EFX_LUT4 LUT__17743 (.I0(n2935), .I1(n7350), .I2(n11538), .O(n7419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17743.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17744 (.I0(n3004), .I1(n7419), .I2(n11596), .O(n7484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17744.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17745 (.I0(n7411), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n7413), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n11601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17745.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17746 (.I0(n2996), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n2998), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n11602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17746.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17747 (.I0(n11602), .I1(n11601), .I2(n11596), .O(n11603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17747.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17748 (.I0(n2933), .I1(n7348), .I2(n11538), .O(n7417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17748.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17749 (.I0(n7415), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n7417), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17749.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17750 (.I0(n11589), .I1(n11567), .I2(n11595), .I3(n11604), 
            .O(n11605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__17750.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__17751 (.I0(n3000), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n3002), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17751.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17752 (.I0(n11567), .I1(n11589), .I2(n11595), .I3(n11606), 
            .O(n11607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__17752.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__17753 (.I0(n11605), .I1(n11607), .O(n11608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__17753.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__17754 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n7484), 
            .I2(n11603), .I3(n11608), .O(n11609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17754.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17755 (.I0(n3000), .I1(n7415), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n11596), .O(n11610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17755.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17756 (.I0(n2998), .I1(n7413), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n11596), .O(n11611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17756.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17757 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n7419), 
            .I2(\u_black_pixel_avg/black_pixel_count[4] ), .I3(n7417), .O(n11612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17757.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17758 (.I0(n11589), .I1(n11567), .I2(n11595), .I3(n11612), 
            .O(n11613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17758.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17759 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n3002), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n3004), .O(n11614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17759.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17760 (.I0(n11567), .I1(n11589), .I2(n11595), .I3(n11614), 
            .O(n11615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__17760.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__17761 (.I0(n11605), .I1(n11607), .I2(n11613), .I3(n11615), 
            .O(n11616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17761.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17762 (.I0(n11611), .I1(n11616), .I2(n11610), .I3(n11603), 
            .O(n11617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__17762.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__17763 (.I0(n2996), .I1(n7411), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11596), .O(n11618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17763.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17764 (.I0(n2994), .I1(n7409), .I2(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I3(n11596), .O(n11619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17764.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17765 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n3240), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n2992), .O(n11620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17765.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17767 (.I0(n11589), .I1(n11620), .I2(n11595), .O(n11622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d3d */ ;
    defparam LUT__17767.LUTMASK = 16'h3d3d;
    EFX_LUT4 LUT__17768 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7655), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7407), .O(n11623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17768.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17769 (.I0(n11567), .I1(n11589), .I2(n11623), .I3(n11595), 
            .O(n11624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__17769.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__17770 (.I0(n11567), .I1(n11622), .I2(n11624), .I3(n11595), 
            .O(n11625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h33e0 */ ;
    defparam LUT__17770.LUTMASK = 16'h33e0;
    EFX_LUT4 LUT__17771 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7651), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n7653), 
            .O(n11626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17771.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17772 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n3236), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n3238), 
            .O(n11627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17772.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17773 (.I0(n11627), .I1(n11626), .I2(n11596), .O(n11628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17773.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17774 (.I0(n11618), .I1(n11619), .I2(n11628), .I3(n11625), 
            .O(n11629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__17774.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__17775 (.I0(n11609), .I1(n11600), .I2(n11617), .I3(n11629), 
            .O(n11630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__17775.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__17776 (.I0(n7407), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n7409), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17776.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17777 (.I0(n2992), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n2994), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17777.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17778 (.I0(n11632), .I1(n11631), .I2(n11596), .O(n11633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17778.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17779 (.I0(n3238), .I1(n7653), .I2(n11596), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17779.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17780 (.I0(n3240), .I1(n7655), .I2(n11596), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17780.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17781 (.I0(n11633), .I1(n11625), .I2(n11634), .I3(n11635), 
            .O(n11636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__17781.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__17782 (.I0(n3275), .I1(n7690), .I2(n11538), .O(n7649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17782.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17783 (.I0(n3234), .I1(n7649), .I2(n11596), .O(n7613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17783.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17784 (.I0(n3236), .I1(n7651), .I2(n11596), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17784.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17785 (.I0(n7645), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n7647), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17785.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17786 (.I0(n3230), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n3232), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17786.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17787 (.I0(n11639), .I1(n11638), .I2(n11596), .O(n11640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17787.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17788 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n7613), 
            .I2(n11637), .I3(n11640), .O(n11641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__17788.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__17789 (.I0(n3228), .I1(n7643), .I2(n11596), .O(n7596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17789.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17790 (.I0(n3226), .I1(n7641), .I2(n11596), .O(n7594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17790.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17791 (.I0(n7594), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n7596), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17791.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17792 (.I0(n11628), .I1(n11636), .I2(n11641), .I3(n11642), 
            .O(n11643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__17792.LUTMASK = 16'he000;
    EFX_LUT4 LUT__17793 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n3222), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n3226), 
            .O(n11644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17793.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17794 (.I0(n3224), .I1(\u_black_pixel_avg/black_pixel_count[18] ), 
            .I2(n11644), .I3(n11596), .O(n11645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h33d0 */ ;
    defparam LUT__17794.LUTMASK = 16'h33d0;
    EFX_LUT4 LUT__17795 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n7641), 
            .I2(\u_black_pixel_avg/black_pixel_count[19] ), .I3(n7637), 
            .O(n11646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17795.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17796 (.I0(n7639), .I1(n11645), .I2(n11646), .I3(n11596), 
            .O(n11647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h70cc */ ;
    defparam LUT__17796.LUTMASK = 16'h70cc;
    EFX_LUT4 LUT__17797 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n7647), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n7649), 
            .O(n11648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17797.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17798 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n3232), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n3234), 
            .O(n11649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17798.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17799 (.I0(n11649), .I1(n11648), .I2(n11596), .O(n11650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17799.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17800 (.I0(n3230), .I1(n7645), .I2(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I3(n11596), .O(n11651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17800.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17801 (.I0(n3228), .I1(n7643), .I2(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I3(n11596), .O(n11652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17801.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17802 (.I0(n11650), .I1(n11640), .I2(n11651), .I3(n11652), 
            .O(n11653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__17802.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__17803 (.I0(n3220), .I1(n7635), .I2(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I3(n11596), .O(n11654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17803.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17804 (.I0(n11567), .I1(n11589), .I2(n11595), .O(n11655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17804.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17805 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n3216), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(n3218), 
            .O(n11656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17805.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17806 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n7631), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(n7633), 
            .O(n11657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17806.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17807 (.I0(n11656), .I1(n11657), .I2(n11655), .O(n11658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17807.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17808 (.I0(n11654), .I1(n11658), .O(n11659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__17808.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__17809 (.I0(n11653), .I1(n11642), .I2(n11647), .I3(n11659), 
            .O(n11660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__17809.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__17810 (.I0(n3222), .I1(n7637), .I2(n11596), .O(n7590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17810.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17811 (.I0(n3224), .I1(n7639), .I2(n11596), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n11661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17811.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17812 (.I0(n7590), .I1(n11661), .I2(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I3(n11654), .O(n11662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__17812.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__17813 (.I0(n3218), .I1(n7633), .I2(n11596), .O(n7586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17813.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17814 (.I0(n3220), .I1(n7635), .I2(n11596), .O(n7588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17814.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17815 (.I0(n7588), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I2(n7586), .I3(\u_black_pixel_avg/black_pixel_count[21] ), 
            .O(n11663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17815.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17816 (.I0(n3255), .I1(n7670), .I2(n11538), .O(n7629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17816.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17817 (.I0(n3214), .I1(n7629), .I2(n11596), .O(n7582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17817.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17818 (.I0(n3216), .I1(n7631), .I2(n11596), .I3(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n11664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17818.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17819 (.I0(n11589), .I1(n11567), .I2(n11595), .I3(n7627), 
            .O(n11665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__17819.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__17820 (.I0(n11567), .I1(n11589), .I2(n11595), .I3(n3212), 
            .O(n11666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__17820.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__17821 (.I0(\u_black_pixel_avg/black_pixel_count[25] ), .I1(n7625), 
            .I2(n10089), .O(n11667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17821.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17822 (.I0(n11666), .I1(n11665), .I2(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I3(n11667), .O(n11668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__17822.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__17823 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(n7582), 
            .I2(n11664), .I3(n11668), .O(n11669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17823.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17824 (.I0(n11662), .I1(n11663), .I2(n11658), .I3(n11669), 
            .O(n11670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__17824.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__17825 (.I0(n11630), .I1(n11643), .I2(n11660), .I3(n11670), 
            .O(n11671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17825.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17826 (.I0(n11665), .I1(n11666), .O(n7580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__17826.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__17827 (.I0(n7580), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[23] ), .I3(n7582), 
            .O(n11672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17827.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17828 (.I0(n3211), .I1(n7625), .I2(n11596), .O(n7578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17828.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17829 (.I0(\u_black_pixel_avg/black_pixel_count[25] ), .I1(n10089), 
            .I2(n7578), .O(n11673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__17829.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__17830 (.I0(n11667), .I1(n11672), .I2(n11673), .O(n11674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__17830.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__17831 (.I0(n11671), .I1(n11674), .O(n11675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17831.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17832 (.I0(n3071), .I1(n7486), .I2(n11675), .O(n7547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17832.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17833 (.I0(\u_black_pixel_avg/y_sum[5] ), .I1(n9702), 
            .O(n11676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17833.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17834 (.I0(n11643), .I1(n11630), .I2(n11660), .O(n11677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__17834.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__17835 (.I0(n11677), .I1(n11670), .I2(n11674), .O(n11678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__17835.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__17836 (.I0(n3075), .I1(\u_black_pixel_avg/y_sum[6] ), 
            .I2(n11676), .I3(n11678), .O(n11679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17836.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17837 (.I0(n3008), .I1(\u_black_pixel_avg/y_sum[7] ), 
            .I2(n11596), .O(n7488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17837.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17838 (.I0(n3073), .I1(n7488), .I2(n11675), .O(n7549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17838.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17839 (.I0(\u_black_pixel_avg/y_sum[5] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17839.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17840 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n7549), 
            .I2(n11679), .I3(n11680), .O(n11681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hddd4 */ ;
    defparam LUT__17840.LUTMASK = 16'hddd4;
    EFX_LUT4 LUT__17841 (.I0(n3071), .I1(n7486), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n11682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17841.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17842 (.I0(n3069), .I1(n7484), .I2(n11675), .O(n7545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17842.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17843 (.I0(n3002), .I1(n7417), .I2(n11596), .O(n7482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17843.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17844 (.I0(n3067), .I1(n7482), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[5] ), 
            .O(n11683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17844.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17845 (.I0(n11682), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n7545), .I3(n11683), .O(n11684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__17845.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__17846 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7484), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n7486), .O(n11685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17846.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17847 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n3069), 
            .I2(\u_black_pixel_avg/black_pixel_count[3] ), .I3(n3071), .O(n11686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17847.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17848 (.I0(n11686), .I1(n11685), .I2(n11675), .O(n11687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17848.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17849 (.I0(n3000), .I1(n7415), .I2(n11596), .O(n7480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17849.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17850 (.I0(n3065), .I1(n7480), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n11675), .O(n11688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17850.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17851 (.I0(n3067), .I1(n7482), .I2(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I3(n11675), .O(n11689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17851.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17852 (.I0(n2994), .I1(n7409), .I2(n11596), .O(n7623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17852.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17853 (.I0(n2992), .I1(n7407), .I2(n11596), .O(n7621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17853.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17854 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7621), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7623), .O(n11690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17854.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17855 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n3207), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n3209), .O(n11691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17855.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17856 (.I0(n11691), .I1(n11690), .I2(n11675), .O(n11692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17856.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17857 (.I0(n2998), .I1(n7413), .I2(n11596), .O(n7478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17857.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17858 (.I0(n2996), .I1(n7411), .I2(n11596), .O(n7476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17858.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17859 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n7476), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n7478), .O(n11693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17859.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17860 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n3061), 
            .I2(\u_black_pixel_avg/black_pixel_count[7] ), .I3(n3063), .O(n11694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17860.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17861 (.I0(n11693), .I1(n11694), .I2(n11671), .I3(n11674), 
            .O(n11695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17861.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17862 (.I0(n11688), .I1(n11689), .I2(n11692), .I3(n11695), 
            .O(n11696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17862.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17863 (.I0(n11681), .I1(n11687), .I2(n11684), .I3(n11696), 
            .O(n11697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__17863.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__17864 (.I0(n7480), .I1(n3065), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__17864.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__17865 (.I0(n7478), .I1(n3063), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[7] ), 
            .O(n11699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__17865.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__17866 (.I0(n3209), .I1(n7623), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[9] ), 
            .O(n11700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17866.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17867 (.I0(n11699), .I1(n11698), .I2(n11695), .I3(n11700), 
            .O(n11701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__17867.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__17868 (.I0(n3061), .I1(n7476), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[8] ), 
            .O(n11702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17868.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17869 (.I0(n3236), .I1(n7651), .I2(n11596), .O(n7615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17869.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17870 (.I0(n3201), .I1(n7615), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[13] ), 
            .O(n11703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17870.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17871 (.I0(n3207), .I1(n7621), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17871.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17872 (.I0(n3240), .I1(n7655), .I2(n11596), .O(n7619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17872.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17873 (.I0(n3205), .I1(n7619), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[11] ), 
            .O(n11705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17873.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17875 (.I0(n3203), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17875.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17876 (.I0(n3238), .I1(n7653), .I2(n11596), .O(n7617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17876.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17877 (.I0(n7617), .I1(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17877.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17878 (.I0(n3232), .I1(n7647), .I2(n11596), .O(n7600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17878.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17879 (.I0(n7600), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n7613), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17879.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17880 (.I0(n3185), .I1(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I2(n3199), .I3(\u_black_pixel_avg/black_pixel_count[14] ), 
            .O(n11710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17880.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17881 (.I0(n11709), .I1(n11710), .I2(n11671), .I3(n11674), 
            .O(n11711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17881.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17882 (.I0(n11707), .I1(n11708), .I2(n11711), .I3(n11678), 
            .O(n11712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17882.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17883 (.I0(n11703), .I1(n11704), .I2(n11705), .I3(n11712), 
            .O(n11713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__17883.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__17884 (.I0(n11702), .I1(n11701), .I2(n11692), .I3(n11713), 
            .O(n11714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__17884.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__17885 (.I0(n3205), .I1(n7619), .I2(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I3(n11675), .O(n11715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17885.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17886 (.I0(n3203), .I1(n7617), .I2(\u_black_pixel_avg/black_pixel_count[12] ), 
            .I3(n11675), .O(n11716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17886.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17887 (.I0(n11716), .I1(n11715), .I2(n11703), .I3(n11712), 
            .O(n11717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__17887.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__17888 (.I0(n3165), .I1(n7580), .I2(\u_black_pixel_avg/black_pixel_count[25] ), 
            .I3(n11675), .O(n11718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17888.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17889 (.I0(n3164), .I1(n7578), .I2(n11675), .I3(n10089), 
            .O(n11719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__17889.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__17890 (.I0(n3167), .I1(n7582), .I2(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I3(n11675), .O(n11720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17890.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17891 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n7588), 
            .I2(\u_black_pixel_avg/black_pixel_count[22] ), .I3(n7586), 
            .O(n11721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17891.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17892 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n3171), 
            .I2(\u_black_pixel_avg/black_pixel_count[21] ), .I3(n3173), 
            .O(n11722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17892.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17893 (.I0(n11721), .I1(n11722), .I2(n11671), .I3(n11674), 
            .O(n11723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17893.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17894 (.I0(n3216), .I1(n7631), .I2(n11596), .O(n7584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17894.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17895 (.I0(n7584), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .I2(n7586), .I3(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n11724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17895.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17896 (.I0(n3169), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .I2(n3171), .I3(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n11725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17896.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17897 (.I0(n11724), .I1(n11725), .I2(n11671), .I3(n11674), 
            .O(n11726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17897.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17898 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(n3169), 
            .O(n11727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17898.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17899 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(n7584), 
            .O(n11728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17899.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17900 (.I0(n11728), .I1(n11727), .I2(n11670), .I3(n11674), 
            .O(n11729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17900.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17901 (.I0(n11727), .I1(n11728), .I2(n11674), .O(n11730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17901.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17902 (.I0(n11730), .I1(n11729), .I2(n11677), .O(n11731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__17902.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__17903 (.I0(n3167), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .O(n11732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17903.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17904 (.I0(n7582), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .O(n11733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17904.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17905 (.I0(n11733), .I1(n11732), .I2(n11670), .I3(n11674), 
            .O(n11734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17905.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17906 (.I0(n11732), .I1(n11733), .I2(n11674), .O(n11735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__17906.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__17907 (.I0(n11735), .I1(n11734), .I2(n11677), .O(n11736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__17907.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__17908 (.I0(n11726), .I1(n11723), .I2(n11731), .I3(n11736), 
            .O(n11737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__17908.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__17909 (.I0(n11718), .I1(n11719), .I2(n11720), .I3(n11737), 
            .O(n11738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17909.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17910 (.I0(n7590), .I1(n3175), .I2(n11671), .I3(n11674), 
            .O(n7537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17910.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17911 (.I0(n3224), .I1(n7639), .I2(n11596), .O(n7592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17911.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17912 (.I0(n7592), .I1(n3177), .I2(n11671), .I3(n11674), 
            .O(n7539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__17912.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__17913 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n7539), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(n7537), 
            .O(n11739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17913.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17914 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n7594), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n7596), 
            .O(n11740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17914.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17915 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n3179), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n3181), 
            .O(n11741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17915.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17916 (.I0(n11740), .I1(n11741), .I2(n11671), .I3(n11674), 
            .O(n11742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__17916.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__17917 (.I0(n11742), .I1(n11739), .O(n11743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17917.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17918 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n7615), 
            .I2(\u_black_pixel_avg/black_pixel_count[14] ), .I3(n7613), 
            .O(n11744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17918.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17919 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n3199), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n3201), 
            .O(n11745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17919.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17920 (.I0(n11745), .I1(n11744), .I2(n11711), .I3(n11675), 
            .O(n11746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17920.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17921 (.I0(n3230), .I1(n7645), .I2(n11596), .O(n7598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17921.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17922 (.I0(n3183), .I1(n7598), .I2(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I3(n11675), .O(n11747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17922.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17923 (.I0(n3185), .I1(n7600), .I2(\u_black_pixel_avg/black_pixel_count[15] ), 
            .I3(n11675), .O(n11748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__17923.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__17924 (.I0(n11746), .I1(n11747), .I2(n11748), .O(n11749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__17924.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__17925 (.I0(n11717), .I1(n11738), .I2(n11743), .I3(n11749), 
            .O(n11750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__17925.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__17926 (.I0(n7594), .I1(n3179), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n11751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__17926.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__17927 (.I0(n7592), .I1(n3177), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n11752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__17927.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__17928 (.I0(n7598), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I2(n7596), .I3(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n11753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17928.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17929 (.I0(n3181), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n3183), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17929.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17930 (.I0(n11754), .I1(n11753), .I2(n11742), .I3(n11675), 
            .O(n11755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__17930.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__17931 (.I0(n11752), .I1(n11751), .I2(n11755), .I3(n11739), 
            .O(n11756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__17931.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__17932 (.I0(n3173), .I1(n7588), .I2(n11675), .O(n7535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17932.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17933 (.I0(n7537), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n11757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17933.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17934 (.I0(n11736), .I1(n11726), .O(n11758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__17934.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__17935 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n7535), 
            .I2(n11757), .I3(n11758), .O(n11759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__17935.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__17936 (.I0(n3164), .I1(n7578), .I2(n11675), .O(n7525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17936.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17937 (.I0(n3165), .I1(n7580), .I2(n11675), .I3(\u_black_pixel_avg/black_pixel_count[25] ), 
            .O(n11760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17937.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17938 (.I0(n7525), .I1(n11760), .I2(\u_black_pixel_avg/black_pixel_count[26] ), 
            .I3(n10490), .O(n11761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b00 */ ;
    defparam LUT__17938.LUTMASK = 16'h2b00;
    EFX_LUT4 LUT__17939 (.I0(n11756), .I1(n11759), .I2(n11738), .I3(n11761), 
            .O(n11762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17939.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17940 (.I0(n11697), .I1(n11714), .I2(n11750), .I3(n11762), 
            .O(n11763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17940.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17941 (.I0(n7547), .I1(n3132), .I2(n11763), .O(n7604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17941.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17942 (.I0(n3199), .I1(n7613), .I2(n11675), .O(n7562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17942.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17943 (.I0(n7562), .I1(n3148), .I2(n11763), .O(n7505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17943.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17944 (.I0(n3185), .I1(n7600), .I2(n11675), .O(n7560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17944.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17945 (.I0(n7560), .I1(n3146), .I2(n11763), .O(n7503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17945.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17946 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n7503), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n7505), 
            .O(n11764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17946.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17947 (.I0(n3203), .I1(n7617), .I2(n11675), .O(n7566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17947.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17948 (.I0(n7566), .I1(n3152), .I2(n11763), .O(n7509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17948.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17949 (.I0(n3201), .I1(n7615), .I2(n11675), .O(n7564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17949.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17950 (.I0(n7564), .I1(n3150), .I2(n11763), .O(n7507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17950.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17951 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n7507), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n7509), 
            .O(n11765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17951.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17952 (.I0(n3205), .I1(n7619), .I2(n11675), .O(n7568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17952.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17953 (.I0(n7568), .I1(n3154), .I2(n11763), .O(n7511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17953.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17954 (.I0(n7509), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n7511), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17954.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17955 (.I0(n7507), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n7505), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n11767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17955.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17956 (.I0(n11766), .I1(n11765), .I2(n11767), .I3(n11764), 
            .O(n11768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__17956.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__17957 (.I0(n3171), .I1(n7586), .I2(n11675), .O(n7533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17957.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17958 (.I0(n7533), .I1(n3118), .I2(n11763), .O(n7474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17958.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17959 (.I0(n7535), .I1(n3120), .I2(n11763), .O(n7491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17959.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17960 (.I0(n7474), .I1(n7491), .I2(\u_black_pixel_avg/black_pixel_count[23] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[22] ), .O(n11769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17960.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17961 (.I0(n3169), .I1(n7584), .I2(n11675), .O(n7531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17961.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17962 (.I0(n7531), .I1(n3116), .I2(n11763), .O(n7472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17962.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17963 (.I0(n3167), .I1(n7582), .I2(n11675), .O(n7529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17963.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17964 (.I0(n7529), .I1(n3114), .I2(n11763), .O(n7470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17964.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17965 (.I0(n7470), .I1(\u_black_pixel_avg/black_pixel_count[25] ), 
            .O(n11770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__17965.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__17966 (.I0(n11769), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I2(n7472), .I3(n11770), .O(n11771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__17966.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__17967 (.I0(n3183), .I1(n7598), .I2(n11675), .O(n7558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17967.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17968 (.I0(n7558), .I1(n3144), .I2(n11763), .O(n7501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17968.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17969 (.I0(n7503), .I1(\u_black_pixel_avg/black_pixel_count[16] ), 
            .I2(n7501), .I3(\u_black_pixel_avg/black_pixel_count[17] ), 
            .O(n11772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17969.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17970 (.I0(n7537), .I1(n3122), .I2(n11763), .I3(\u_black_pixel_avg/black_pixel_count[21] ), 
            .O(n11773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17970.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17971 (.I0(n7539), .I1(n3124), .I2(n11763), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n11774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17971.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17972 (.I0(n3179), .I1(n7594), .I2(n11675), .O(n7554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17972.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17973 (.I0(n7554), .I1(n3140), .I2(n11763), .I3(\u_black_pixel_avg/black_pixel_count[19] ), 
            .O(n11775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17973.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17974 (.I0(n3181), .I1(n7596), .I2(n11675), .O(n7556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17974.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17975 (.I0(n7556), .I1(n3142), .I2(n11763), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n11776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__17975.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__17976 (.I0(n11773), .I1(n11774), .I2(n11775), .I3(n11776), 
            .O(n11777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__17976.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__17977 (.I0(n11768), .I1(n11771), .I2(n11772), .I3(n11777), 
            .O(n11778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__17977.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__17978 (.I0(n3075), .I1(\u_black_pixel_avg/y_sum[6] ), 
            .I2(n11675), .O(n7551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17978.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17979 (.I0(\u_black_pixel_avg/y_sum[5] ), .I1(\u_black_pixel_avg/y_sum[4] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__17979.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__17980 (.I0(n7551), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n11779), .O(n11780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__17980.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__17981 (.I0(n7549), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n11763), .I3(n11780), .O(n11781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__17981.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__17982 (.I0(n7549), .I1(n3134), .I2(n11763), .O(n7606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17982.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17983 (.I0(n7606), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n11781), .O(n11782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__17983.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__17984 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n3138), 
            .I2(\u_black_pixel_avg/y_sum[4] ), .I3(\u_black_pixel_avg/black_pixel_count[0] ), 
            .O(n11783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__17984.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__17985 (.I0(n11783), .I1(n3136), .I2(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n11784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__17985.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__17986 (.I0(n3134), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(n11784), .O(n11785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__17986.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__17987 (.I0(n11763), .I1(n11785), .I2(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I3(n7604), .O(n11786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__17987.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__17988 (.I0(n7545), .I1(n3130), .I2(n11763), .O(n7602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17988.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17989 (.I0(n7602), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n7604), .I3(\u_black_pixel_avg/black_pixel_count[4] ), .O(n11787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17989.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17990 (.I0(n3067), .I1(n7482), .I2(n11675), .O(n7543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17990.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17991 (.I0(n7543), .I1(n3128), .I2(n11763), .O(n7523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17991.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17992 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n7523), 
            .I2(\u_black_pixel_avg/black_pixel_count[5] ), .I3(n7602), .O(n11788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17992.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17993 (.I0(n11786), .I1(n11782), .I2(n11787), .I3(n11788), 
            .O(n11789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__17993.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__17994 (.I0(n3063), .I1(n7478), .I2(n11675), .O(n7576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17994.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17995 (.I0(n7576), .I1(n3162), .I2(n11763), .O(n7519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17995.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17996 (.I0(n3061), .I1(n7476), .I2(n11675), .O(n7574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17996.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17997 (.I0(n7574), .I1(n3160), .I2(n11763), .O(n7517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17997.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__17998 (.I0(n7517), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n7519), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__17998.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__17999 (.I0(n3065), .I1(n7480), .I2(n11675), .O(n7541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__17999.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18000 (.I0(n7541), .I1(n3126), .I2(n11763), .O(n7521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18000.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18001 (.I0(n7521), .I1(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I2(n7523), .I3(\u_black_pixel_avg/black_pixel_count[6] ), .O(n11791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18001.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18002 (.I0(n3209), .I1(n7623), .I2(n11675), .O(n7572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18002.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18003 (.I0(n7572), .I1(n3158), .I2(n11763), .O(n7515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18003.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18004 (.I0(n3207), .I1(n7621), .I2(n11675), .O(n7570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18004.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18005 (.I0(n7570), .I1(n3156), .I2(n11763), .O(n7513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18005.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18006 (.I0(n7513), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n7515), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18006.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18007 (.I0(n11790), .I1(n11791), .I2(n11792), .O(n11793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18007.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18008 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n7521), 
            .I2(\u_black_pixel_avg/black_pixel_count[8] ), .I3(n7519), .O(n11794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18008.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18009 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n7515), 
            .I2(\u_black_pixel_avg/black_pixel_count[9] ), .I3(n7517), .O(n11795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18009.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18010 (.I0(n11794), .I1(n11790), .I2(n11795), .I3(n11792), 
            .O(n11796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__18010.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__18011 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7511), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n7513), 
            .O(n11797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18011.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18012 (.I0(n11797), .I1(n11764), .I2(n11765), .O(n11798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18012.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18013 (.I0(n11793), .I1(n11789), .I2(n11796), .I3(n11798), 
            .O(n11799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__18013.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__18014 (.I0(n7525), .I1(n3111), .I2(n11763), .O(n7466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18014.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18015 (.I0(n3165), .I1(n7580), .I2(n11675), .O(n7527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18015.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18016 (.I0(n7527), .I1(n3112), .I2(n11763), .O(n7468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18016.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18017 (.I0(n7466), .I1(n7468), .I2(\u_black_pixel_avg/black_pixel_count[27] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[26] ), .O(n11800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__18017.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__18018 (.I0(\u_black_pixel_avg/black_pixel_count[28] ), .I1(n10489), 
            .I2(n11800), .O(n11801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__18018.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__18019 (.I0(n7556), .I1(n3142), .I2(n11763), .O(n7499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18019.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18020 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n7501), 
            .I2(\u_black_pixel_avg/black_pixel_count[18] ), .I3(n7499), 
            .O(n11802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18020.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18021 (.I0(n11802), .I1(n11777), .O(n11803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18021.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18022 (.I0(n7539), .I1(n3124), .I2(n11763), .O(n7495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18022.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18023 (.I0(n7554), .I1(n3140), .I2(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I3(n11763), .O(n11804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__18023.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__18024 (.I0(n7495), .I1(\u_black_pixel_avg/black_pixel_count[20] ), 
            .I2(n11804), .I3(n11773), .O(n11805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__18024.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__18025 (.I0(\u_black_pixel_avg/black_pixel_count[24] ), .I1(n7472), 
            .I2(\u_black_pixel_avg/black_pixel_count[23] ), .I3(n7474), 
            .O(n11806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18025.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18026 (.I0(n7537), .I1(n3122), .I2(n11763), .O(n7493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18026.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18027 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n7493), 
            .I2(\u_black_pixel_avg/black_pixel_count[22] ), .I3(n7491), 
            .O(n11807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18027.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18028 (.I0(n11805), .I1(n11806), .I2(n11807), .O(n11808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__18028.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__18029 (.I0(\u_black_pixel_avg/black_pixel_count[25] ), .I1(n7470), 
            .I2(\u_black_pixel_avg/black_pixel_count[27] ), .I3(n7466), 
            .O(n11809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18029.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18030 (.I0(\u_black_pixel_avg/black_pixel_count[26] ), .I1(n7468), 
            .I2(n11809), .O(n11810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__18030.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__18031 (.I0(n11803), .I1(n11808), .I2(n11771), .I3(n11810), 
            .O(n11811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__18031.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__18032 (.I0(n11799), .I1(n11778), .I2(n11811), .I3(n11801), 
            .O(n11812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__18032.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__18033 (.I0(n3189), .I1(n7604), .I2(n11812), .O(n7464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18033.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18034 (.I0(n3191), .I1(n7606), .I2(n11812), .I3(\u_black_pixel_avg/black_pixel_count[4] ), 
            .O(n11813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__18034.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__18035 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n7464), 
            .I2(n11813), .O(n11814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__18035.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__18036 (.I0(\u_black_pixel_avg/y_sum[3] ), .I1(\u_black_pixel_avg/black_pixel_count[0] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[1] ), .O(n11815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__18036.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__18037 (.I0(n3197), .I1(\u_black_pixel_avg/y_sum[4] ), 
            .I2(n11815), .I3(n11812), .O(n11816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__18037.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__18038 (.I0(\u_black_pixel_avg/y_sum[5] ), .I1(n3138), 
            .I2(n11763), .O(n7610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18038.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18039 (.I0(n3195), .I1(n7610), .I2(n11812), .I3(\u_black_pixel_avg/black_pixel_count[2] ), 
            .O(n11817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__18039.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__18040 (.I0(n7551), .I1(n3136), .I2(n11763), .O(n7608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18040.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18041 (.I0(n3193), .I1(n7608), .I2(n11812), .I3(\u_black_pixel_avg/black_pixel_count[3] ), 
            .O(n11818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__18041.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__18042 (.I0(\u_black_pixel_avg/y_sum[3] ), .I1(n9702), 
            .O(n11819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18042.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18043 (.I0(n11816), .I1(n11817), .I2(n11818), .I3(n11819), 
            .O(n11820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__18043.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__18044 (.I0(n7608), .I1(\u_black_pixel_avg/black_pixel_count[3] ), 
            .I2(\u_black_pixel_avg/black_pixel_count[2] ), .I3(n7610), .O(n11821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__18044.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__18045 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n7606), 
            .I2(n11821), .O(n11822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__18045.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__18046 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(\u_black_pixel_avg/black_pixel_count[2] ), 
            .I2(n3193), .I3(n3195), .O(n11823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__18046.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__18047 (.I0(n3191), .I1(\u_black_pixel_avg/black_pixel_count[4] ), 
            .I2(n11823), .O(n11824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__18047.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__18048 (.I0(n11824), .I1(n11822), .I2(n11812), .O(n11825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18048.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18049 (.I0(n7464), .I1(\u_black_pixel_avg/black_pixel_count[5] ), 
            .I2(n11813), .I3(n11825), .O(n11826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hddd4 */ ;
    defparam LUT__18049.LUTMASK = 16'hddd4;
    EFX_LUT4 LUT__18050 (.I0(n3109), .I1(n7523), .I2(n11812), .O(n7460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18050.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18051 (.I0(n3187), .I1(n7602), .I2(\u_black_pixel_avg/black_pixel_count[6] ), 
            .I3(n11812), .O(n11827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__18051.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__18052 (.I0(n3107), .I1(n7521), .I2(\u_black_pixel_avg/black_pixel_count[8] ), 
            .I3(n11812), .O(n11828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__18052.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__18053 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n7460), 
            .I2(n11827), .I3(n11828), .O(n11829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__18053.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__18054 (.I0(n11820), .I1(n11814), .I2(n11826), .I3(n11829), 
            .O(n11830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__18054.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__18055 (.I0(n3187), .I1(n7602), .I2(n11812), .I3(\u_black_pixel_avg/black_pixel_count[6] ), 
            .O(n11831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__18055.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__18056 (.I0(n7460), .I1(n11831), .I2(\u_black_pixel_avg/black_pixel_count[7] ), 
            .I3(n11828), .O(n11832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__18056.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__18057 (.I0(n3103), .I1(n7517), .I2(n11812), .O(n7454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18057.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18058 (.I0(n3101), .I1(n7515), .I2(n11812), .O(n7452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18058.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18059 (.I0(n7452), .I1(\u_black_pixel_avg/black_pixel_count[11] ), 
            .I2(n7454), .I3(\u_black_pixel_avg/black_pixel_count[10] ), 
            .O(n11833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18059.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18060 (.I0(n3099), .I1(n7513), .I2(n11812), .O(n7450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18060.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18061 (.I0(n3097), .I1(n7511), .I2(n11812), .O(n7448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18061.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18062 (.I0(n7448), .I1(\u_black_pixel_avg/black_pixel_count[13] ), 
            .I2(n7450), .I3(\u_black_pixel_avg/black_pixel_count[12] ), 
            .O(n11834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18062.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18063 (.I0(n3107), .I1(n7521), .I2(n11812), .O(n7458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18063.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18064 (.I0(n3105), .I1(n7519), .I2(n11812), .O(n7456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18064.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18065 (.I0(n7456), .I1(\u_black_pixel_avg/black_pixel_count[9] ), 
            .I2(n7458), .I3(\u_black_pixel_avg/black_pixel_count[8] ), .O(n11835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18065.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18066 (.I0(n11832), .I1(n11833), .I2(n11834), .I3(n11835), 
            .O(n11836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__18066.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__18067 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n7456), 
            .I2(\u_black_pixel_avg/black_pixel_count[10] ), .I3(n7454), 
            .O(n11837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18067.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18068 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n7450), 
            .I2(\u_black_pixel_avg/black_pixel_count[11] ), .I3(n7452), 
            .O(n11838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18068.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18069 (.I0(n11837), .I1(n11833), .I2(n11838), .I3(n11834), 
            .O(n11839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__18069.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__18070 (.I0(n3093), .I1(n7507), .I2(n11812), .O(n7444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18070.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18071 (.I0(n3091), .I1(n7505), .I2(n11812), .O(n7442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18071.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18072 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n7442), 
            .I2(\u_black_pixel_avg/black_pixel_count[15] ), .I3(n7444), 
            .O(n11840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18072.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18073 (.I0(n3095), .I1(n7509), .I2(n11812), .O(n7446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18073.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18074 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n7446), 
            .I2(\u_black_pixel_avg/black_pixel_count[13] ), .I3(n7448), 
            .O(n11841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18074.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18075 (.I0(n3089), .I1(n7503), .I2(n11812), .O(n7440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18075.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18076 (.I0(n3087), .I1(n7501), .I2(n11812), .O(n7438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18076.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18077 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n7438), 
            .I2(\u_black_pixel_avg/black_pixel_count[17] ), .I3(n7440), 
            .O(n11842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18077.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18078 (.I0(n11840), .I1(n11841), .I2(n11842), .O(n11843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18078.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18079 (.I0(n11836), .I1(n11830), .I2(n11839), .I3(n11843), 
            .O(n11844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__18079.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__18080 (.I0(n7446), .I1(\u_black_pixel_avg/black_pixel_count[14] ), 
            .I2(n7444), .I3(\u_black_pixel_avg/black_pixel_count[15] ), 
            .O(n11845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18080.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18081 (.I0(n7440), .I1(\u_black_pixel_avg/black_pixel_count[17] ), 
            .I2(n7442), .I3(\u_black_pixel_avg/black_pixel_count[16] ), 
            .O(n11846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18081.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18082 (.I0(n11845), .I1(n11840), .I2(n11846), .I3(n11842), 
            .O(n11847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__18082.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__18083 (.I0(n3079), .I1(n7493), .I2(n11812), .O(n7430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18083.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18084 (.I0(n3077), .I1(n7491), .I2(n11812), .O(n7428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18084.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18085 (.I0(n7428), .I1(\u_black_pixel_avg/black_pixel_count[23] ), 
            .I2(n7430), .I3(\u_black_pixel_avg/black_pixel_count[22] ), 
            .O(n11848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18085.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18086 (.I0(n7554), .I1(n3140), .I2(n11763), .O(n7497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18086.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18087 (.I0(n3083), .I1(n7497), .I2(n11812), .O(n7434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18087.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18088 (.I0(n3081), .I1(n7495), .I2(n11812), .O(n7432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18088.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18089 (.I0(n7432), .I1(\u_black_pixel_avg/black_pixel_count[21] ), 
            .I2(n7434), .I3(\u_black_pixel_avg/black_pixel_count[20] ), 
            .O(n11849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18089.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18090 (.I0(n3085), .I1(n7499), .I2(n11812), .O(n7436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18090.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18091 (.I0(n7436), .I1(\u_black_pixel_avg/black_pixel_count[19] ), 
            .I2(n7438), .I3(\u_black_pixel_avg/black_pixel_count[18] ), 
            .O(n11850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18091.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18092 (.I0(n11847), .I1(n11848), .I2(n11849), .I3(n11850), 
            .O(n11851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__18092.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__18093 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n7436), 
            .I2(\u_black_pixel_avg/black_pixel_count[20] ), .I3(n7434), 
            .O(n11852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18093.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18094 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n7432), 
            .I2(\u_black_pixel_avg/black_pixel_count[22] ), .I3(n7430), 
            .O(n11853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18094.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18095 (.I0(n11852), .I1(n11849), .I2(n11853), .I3(n11848), 
            .O(n11854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__18095.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__18096 (.I0(n3055), .I1(n7470), .I2(n11812), .O(n7405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18096.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18097 (.I0(n3052), .I1(n7466), .I2(n11812), .O(n7401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18097.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18098 (.I0(\u_black_pixel_avg/black_pixel_count[28] ), .I1(n7401), 
            .O(n11855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18098.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18099 (.I0(n3053), .I1(n7468), .I2(n11812), .O(n7403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18099.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18100 (.I0(n3057), .I1(n7472), .I2(n11812), .O(n7424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18100.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18101 (.I0(\u_black_pixel_avg/black_pixel_count[25] ), .I1(n7424), 
            .I2(\u_black_pixel_avg/black_pixel_count[27] ), .I3(n7403), 
            .O(n11856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18101.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18102 (.I0(\u_black_pixel_avg/black_pixel_count[26] ), .I1(n7405), 
            .I2(n11855), .I3(n11856), .O(n11857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__18102.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__18103 (.I0(n3059), .I1(n7474), .I2(n11812), .O(n7426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18103.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18104 (.I0(\u_black_pixel_avg/black_pixel_count[24] ), .I1(n7426), 
            .I2(\u_black_pixel_avg/black_pixel_count[23] ), .I3(n7428), 
            .O(n11858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18104.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18105 (.I0(n11854), .I1(n11857), .I2(n11858), .O(n11859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__18105.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__18106 (.I0(n7426), .I1(\u_black_pixel_avg/black_pixel_count[24] ), 
            .I2(n7424), .I3(\u_black_pixel_avg/black_pixel_count[25] ), 
            .O(n11860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__18106.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__18107 (.I0(n7403), .I1(n7405), .I2(\u_black_pixel_avg/black_pixel_count[27] ), 
            .I3(\u_black_pixel_avg/black_pixel_count[26] ), .O(n11861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__18107.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__18108 (.I0(n11855), .I1(n11861), .O(n11862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__18108.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__18109 (.I0(\u_black_pixel_avg/black_pixel_count[28] ), .I1(n7466), 
            .I2(n10489), .O(n11863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__18109.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__18110 (.I0(n11860), .I1(n11857), .I2(n11862), .I3(n11863), 
            .O(n11864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__18110.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__18111 (.I0(n11844), .I1(n11851), .I2(n11859), .I3(n11864), 
            .O(n11865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__18111.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__18391 (.I0(\u_black_pixel_avg/x_sum[1] ), .I1(n4074), 
            .I2(n9701), .O(\u_black_pixel_avg/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18391.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18392 (.I0(\u_black_pixel_avg/x_sum[0] ), .I1(n1714), 
            .I2(n9701), .O(\u_black_pixel_avg/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18392.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18393 (.I0(\u_black_pixel_avg/y_sum[1] ), .I1(n4013), 
            .I2(n9701), .O(\u_black_pixel_avg/n174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18393.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18394 (.I0(\u_black_pixel_avg/y_sum[2] ), .I1(n4011), 
            .I2(n9701), .O(\u_black_pixel_avg/n173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18394.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18395 (.I0(\u_black_pixel_avg/y_sum[3] ), .I1(n4009), 
            .I2(n9701), .O(\u_black_pixel_avg/n172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18395.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18396 (.I0(\u_black_pixel_avg/y_sum[4] ), .I1(n4007), 
            .I2(n9701), .O(\u_black_pixel_avg/n171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18396.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18397 (.I0(\u_black_pixel_avg/y_sum[5] ), .I1(n4005), 
            .I2(n9701), .O(\u_black_pixel_avg/n170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18397.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18398 (.I0(\u_black_pixel_avg/y_sum[6] ), .I1(n4003), 
            .I2(n9701), .O(\u_black_pixel_avg/n169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18398.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18399 (.I0(\u_black_pixel_avg/y_sum[7] ), .I1(n4001), 
            .I2(n9701), .O(\u_black_pixel_avg/n168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18399.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18400 (.I0(\u_black_pixel_avg/y_sum[8] ), .I1(n3999), 
            .I2(n9701), .O(\u_black_pixel_avg/n167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18400.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18401 (.I0(\u_black_pixel_avg/y_sum[9] ), .I1(n3997), 
            .I2(n9701), .O(\u_black_pixel_avg/n166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18401.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18402 (.I0(\u_black_pixel_avg/y_sum[10] ), .I1(n3995), 
            .I2(n9701), .O(\u_black_pixel_avg/n165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18402.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18403 (.I0(\u_black_pixel_avg/y_sum[11] ), .I1(n3993), 
            .I2(n9701), .O(\u_black_pixel_avg/n164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18403.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18404 (.I0(\u_black_pixel_avg/y_sum[12] ), .I1(n3991), 
            .I2(n9701), .O(\u_black_pixel_avg/n163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18404.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18405 (.I0(\u_black_pixel_avg/y_sum[13] ), .I1(n3989), 
            .I2(n9701), .O(\u_black_pixel_avg/n162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18405.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18406 (.I0(\u_black_pixel_avg/y_sum[14] ), .I1(n3987), 
            .I2(n9701), .O(\u_black_pixel_avg/n161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18406.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18407 (.I0(\u_black_pixel_avg/y_sum[15] ), .I1(n3985), 
            .I2(n9701), .O(\u_black_pixel_avg/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18407.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18408 (.I0(\u_black_pixel_avg/y_sum[16] ), .I1(n3983), 
            .I2(n9701), .O(\u_black_pixel_avg/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18408.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18409 (.I0(\u_black_pixel_avg/y_sum[17] ), .I1(n3981), 
            .I2(n9701), .O(\u_black_pixel_avg/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18409.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18410 (.I0(\u_black_pixel_avg/y_sum[18] ), .I1(n3979), 
            .I2(n9701), .O(\u_black_pixel_avg/n157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18410.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18411 (.I0(\u_black_pixel_avg/y_sum[19] ), .I1(n3977), 
            .I2(n9701), .O(\u_black_pixel_avg/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18411.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18412 (.I0(\u_black_pixel_avg/y_sum[20] ), .I1(n3975), 
            .I2(n9701), .O(\u_black_pixel_avg/n155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18412.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18413 (.I0(\u_black_pixel_avg/y_sum[21] ), .I1(n3973), 
            .I2(n9701), .O(\u_black_pixel_avg/n154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18413.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18414 (.I0(\u_black_pixel_avg/y_sum[22] ), .I1(n3971), 
            .I2(n9701), .O(\u_black_pixel_avg/n153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18414.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18415 (.I0(\u_black_pixel_avg/y_sum[23] ), .I1(n3969), 
            .I2(n9701), .O(\u_black_pixel_avg/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18415.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18416 (.I0(\u_black_pixel_avg/y_sum[24] ), .I1(n3967), 
            .I2(n9701), .O(\u_black_pixel_avg/n151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18416.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18417 (.I0(\u_black_pixel_avg/y_sum[25] ), .I1(n3965), 
            .I2(n9701), .O(\u_black_pixel_avg/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18417.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18418 (.I0(\u_black_pixel_avg/y_sum[26] ), .I1(n3963), 
            .I2(n9701), .O(\u_black_pixel_avg/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18418.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18419 (.I0(\u_black_pixel_avg/y_sum[27] ), .I1(n3961), 
            .I2(n9701), .O(\u_black_pixel_avg/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18419.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18420 (.I0(\u_black_pixel_avg/y_sum[28] ), .I1(n3959), 
            .I2(n9701), .O(\u_black_pixel_avg/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18420.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18421 (.I0(\u_black_pixel_avg/y_sum[29] ), .I1(n3957), 
            .I2(n9701), .O(\u_black_pixel_avg/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18421.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18422 (.I0(\u_black_pixel_avg/y_sum[30] ), .I1(n3955), 
            .I2(n9701), .O(\u_black_pixel_avg/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18422.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18423 (.I0(\u_black_pixel_avg/y_sum[31] ), .I1(n3954), 
            .I2(n9701), .O(\u_black_pixel_avg/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18423.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18424 (.I0(\u_black_pixel_avg/black_pixel_count[1] ), .I1(n1679), 
            .I2(n9701), .O(\u_black_pixel_avg/n207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18424.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18425 (.I0(\u_black_pixel_avg/black_pixel_count[2] ), .I1(n4133), 
            .I2(n9701), .O(\u_black_pixel_avg/n206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18425.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18426 (.I0(\u_black_pixel_avg/black_pixel_count[3] ), .I1(n4131), 
            .I2(n9701), .O(\u_black_pixel_avg/n205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18426.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18427 (.I0(\u_black_pixel_avg/black_pixel_count[4] ), .I1(n4129), 
            .I2(n9701), .O(\u_black_pixel_avg/n204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18427.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18428 (.I0(\u_black_pixel_avg/black_pixel_count[5] ), .I1(n4127), 
            .I2(n9701), .O(\u_black_pixel_avg/n203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18428.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18429 (.I0(\u_black_pixel_avg/black_pixel_count[6] ), .I1(n4125), 
            .I2(n9701), .O(\u_black_pixel_avg/n202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18429.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18430 (.I0(\u_black_pixel_avg/black_pixel_count[7] ), .I1(n4123), 
            .I2(n9701), .O(\u_black_pixel_avg/n201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18430.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18431 (.I0(\u_black_pixel_avg/black_pixel_count[8] ), .I1(n4121), 
            .I2(n9701), .O(\u_black_pixel_avg/n200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18431.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18432 (.I0(\u_black_pixel_avg/black_pixel_count[9] ), .I1(n4119), 
            .I2(n9701), .O(\u_black_pixel_avg/n199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18432.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18433 (.I0(\u_black_pixel_avg/black_pixel_count[10] ), .I1(n4117), 
            .I2(n9701), .O(\u_black_pixel_avg/n198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18433.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18434 (.I0(\u_black_pixel_avg/black_pixel_count[11] ), .I1(n4115), 
            .I2(n9701), .O(\u_black_pixel_avg/n197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18434.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18435 (.I0(\u_black_pixel_avg/black_pixel_count[12] ), .I1(n4113), 
            .I2(n9701), .O(\u_black_pixel_avg/n196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18435.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18436 (.I0(\u_black_pixel_avg/black_pixel_count[13] ), .I1(n4111), 
            .I2(n9701), .O(\u_black_pixel_avg/n195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18436.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18437 (.I0(\u_black_pixel_avg/black_pixel_count[14] ), .I1(n4109), 
            .I2(n9701), .O(\u_black_pixel_avg/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18437.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18438 (.I0(\u_black_pixel_avg/black_pixel_count[15] ), .I1(n4107), 
            .I2(n9701), .O(\u_black_pixel_avg/n193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18438.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18439 (.I0(\u_black_pixel_avg/black_pixel_count[16] ), .I1(n4105), 
            .I2(n9701), .O(\u_black_pixel_avg/n192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18439.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18440 (.I0(\u_black_pixel_avg/black_pixel_count[17] ), .I1(n4103), 
            .I2(n9701), .O(\u_black_pixel_avg/n191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18440.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18441 (.I0(\u_black_pixel_avg/black_pixel_count[18] ), .I1(n4101), 
            .I2(n9701), .O(\u_black_pixel_avg/n190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18441.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18442 (.I0(\u_black_pixel_avg/black_pixel_count[19] ), .I1(n4099), 
            .I2(n9701), .O(\u_black_pixel_avg/n189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18442.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18443 (.I0(\u_black_pixel_avg/black_pixel_count[20] ), .I1(n4097), 
            .I2(n9701), .O(\u_black_pixel_avg/n188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18443.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18444 (.I0(\u_black_pixel_avg/black_pixel_count[21] ), .I1(n4095), 
            .I2(n9701), .O(\u_black_pixel_avg/n187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18444.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18445 (.I0(\u_black_pixel_avg/black_pixel_count[22] ), .I1(n4093), 
            .I2(n9701), .O(\u_black_pixel_avg/n186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18445.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18446 (.I0(\u_black_pixel_avg/black_pixel_count[23] ), .I1(n4091), 
            .I2(n9701), .O(\u_black_pixel_avg/n185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18446.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18447 (.I0(\u_black_pixel_avg/black_pixel_count[24] ), .I1(n4089), 
            .I2(n9701), .O(\u_black_pixel_avg/n184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18447.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18448 (.I0(\u_black_pixel_avg/black_pixel_count[25] ), .I1(n4087), 
            .I2(n9701), .O(\u_black_pixel_avg/n183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18448.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18449 (.I0(\u_black_pixel_avg/black_pixel_count[26] ), .I1(n4085), 
            .I2(n9701), .O(\u_black_pixel_avg/n182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18449.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18450 (.I0(\u_black_pixel_avg/black_pixel_count[27] ), .I1(n4083), 
            .I2(n9701), .O(\u_black_pixel_avg/n181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18450.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18451 (.I0(\u_black_pixel_avg/black_pixel_count[28] ), .I1(n4081), 
            .I2(n9701), .O(\u_black_pixel_avg/n180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18451.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18452 (.I0(\u_black_pixel_avg/black_pixel_count[29] ), .I1(n4079), 
            .I2(n9701), .O(\u_black_pixel_avg/n179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18452.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18453 (.I0(\u_black_pixel_avg/black_pixel_count[30] ), .I1(n4077), 
            .I2(n9701), .O(\u_black_pixel_avg/n178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18453.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18454 (.I0(\u_black_pixel_avg/black_pixel_count[31] ), .I1(n4076), 
            .I2(n9701), .O(\u_black_pixel_avg/n177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18454.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18460 (.I0(\x_avg_black[6] ), .I1(n10455), .I2(n10838), 
            .O(\u_black_pixel_avg/n483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18460.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18461 (.I0(\x_avg_black[7] ), .I1(n10400), .I2(n10838), 
            .O(\u_black_pixel_avg/n482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18461.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18462 (.I0(\x_avg_black[8] ), .I1(n10336), .I2(n10838), 
            .O(\u_black_pixel_avg/n481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18462.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18463 (.I0(\x_avg_black[9] ), .I1(n10293), .I2(n10838), 
            .O(\u_black_pixel_avg/n480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18463.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18464 (.I0(\x_avg_black[10] ), .I1(n10255), .I2(n10838), 
            .O(\u_black_pixel_avg/n479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18464.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18465 (.I0(\x_avg_black[11] ), .I1(n10215), .I2(n10838), 
            .O(\u_black_pixel_avg/n478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18465.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18466 (.I0(n9734), .I1(n9735), .O(n6202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__18466.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__18467 (.I0(n10856), .I1(n10864), .O(n6759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__18467.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__18468 (.I0(\u_lcd_driver/r_lcd_dv ), .I1(\u_lcd_driver/r_lcd_rgb[23] ), 
            .O(n7221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18468.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18469 (.I0(n7221), .I1(\u_rgb2dvi/enc_2/acc[4] ), .O(\u_rgb2dvi/enc_2/q_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18469.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18470 (.I0(n2812), .I1(n2838), .I2(\u_rgb2dvi/enc_2/q_out[9] ), 
            .O(n12080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18470.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18471 (.I0(n2824), .I1(n2817), .I2(n7221), .O(n12081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18471.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18472 (.I0(\u_rgb2dvi/enc_2/acc[0] ), .I1(\u_rgb2dvi/enc_2/acc[1] ), 
            .I2(\u_rgb2dvi/enc_2/acc[2] ), .I3(\u_rgb2dvi/enc_2/acc[3] ), 
            .O(n12082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__18472.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__18473 (.I0(\u_rgb2dvi/enc_2/acc[4] ), .I1(n12082), .O(n12083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18473.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18474 (.I0(n12081), .I1(n12080), .I2(n12083), .O(n7160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18474.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18475 (.I0(n2813), .I1(n2779), .I2(\u_rgb2dvi/enc_2/q_out[9] ), 
            .O(n12084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18475.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18476 (.I0(n2825), .I1(n2818), .I2(n7221), .O(n12085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18476.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18477 (.I0(n12085), .I1(n12084), .I2(n12083), .O(n7163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18477.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18478 (.I0(n2815), .I1(n3350), .I2(\u_rgb2dvi/enc_2/q_out[9] ), 
            .O(n12086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18478.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18479 (.I0(n2827), .I1(n2820), .I2(n7221), .O(n12087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18479.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18480 (.I0(n12087), .I1(n12086), .I2(n12083), .O(n7166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18480.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18481 (.I0(n3468), .I1(n3352), .I2(\u_rgb2dvi/enc_2/q_out[9] ), 
            .O(n12088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18481.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18482 (.I0(n2829), .I1(n2822), .I2(n7221), .O(n12089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18482.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18483 (.I0(n12089), .I1(n12088), .I2(n12083), .O(n7169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18483.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18484 (.I0(n7221), .I1(\u_rgb2dvi/enc_1/acc[4] ), .O(\u_rgb2dvi/enc_1/q_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18484.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18485 (.I0(n2812), .I1(n2838), .I2(\u_rgb2dvi/enc_1/q_out[9] ), 
            .O(n12090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18485.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18486 (.I0(\u_rgb2dvi/enc_1/acc[0] ), .I1(\u_rgb2dvi/enc_1/acc[1] ), 
            .I2(\u_rgb2dvi/enc_1/acc[2] ), .I3(\u_rgb2dvi/enc_1/acc[3] ), 
            .O(n12091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__18486.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__18487 (.I0(\u_rgb2dvi/enc_1/acc[4] ), .I1(n12091), .O(n12092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18487.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18488 (.I0(n12081), .I1(n12090), .I2(n12092), .O(n7174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18488.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18489 (.I0(n2813), .I1(n2779), .I2(\u_rgb2dvi/enc_1/q_out[9] ), 
            .O(n12093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18489.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18490 (.I0(n12085), .I1(n12093), .I2(n12092), .O(n7177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18490.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18491 (.I0(n2815), .I1(n3350), .I2(\u_rgb2dvi/enc_1/q_out[9] ), 
            .O(n12094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18491.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18492 (.I0(n12087), .I1(n12094), .I2(n12092), .O(n7180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18492.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18493 (.I0(n3468), .I1(n3352), .I2(\u_rgb2dvi/enc_1/q_out[9] ), 
            .O(n12095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18493.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18494 (.I0(n12089), .I1(n12095), .I2(n12092), .O(n7183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18494.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18495 (.I0(n2812), .I1(n2838), .I2(n7221), .I3(\u_rgb2dvi/enc_0/acc[4] ), 
            .O(n12096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__18495.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__18496 (.I0(\u_rgb2dvi/enc_0/acc[0] ), .I1(\u_rgb2dvi/enc_0/acc[1] ), 
            .I2(\u_rgb2dvi/enc_0/acc[2] ), .I3(\u_rgb2dvi/enc_0/acc[3] ), 
            .O(n12097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__18496.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__18497 (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(n12097), .O(n12098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18497.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18498 (.I0(n12096), .I1(n12081), .I2(n12098), .O(n7226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18498.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18499 (.I0(n2779), .I1(n2813), .I2(n7221), .I3(\u_rgb2dvi/enc_0/acc[4] ), 
            .O(n12099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__18499.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__18500 (.I0(n12099), .I1(n12085), .I2(n12098), .O(n7229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18500.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18501 (.I0(n2815), .I1(n3350), .I2(n7221), .I3(\u_rgb2dvi/enc_0/acc[4] ), 
            .O(n12100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__18501.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__18502 (.I0(n12100), .I1(n12087), .I2(n12098), .O(n7232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18502.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18503 (.I0(n3352), .I1(n3468), .I2(n7221), .I3(\u_rgb2dvi/enc_0/acc[4] ), 
            .O(n12101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__18503.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__18504 (.I0(n12101), .I1(n12089), .I2(n12098), .O(n7235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18504.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18507 (.I0(\y_avg_black[3] ), .I1(n11865), .I2(n10838), 
            .O(\u_black_pixel_avg/n499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18507.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18508 (.I0(\y_avg_black[4] ), .I1(n11812), .I2(n10838), 
            .O(\u_black_pixel_avg/n498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18508.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18509 (.I0(\y_avg_black[5] ), .I1(n11763), .I2(n10838), 
            .O(\u_black_pixel_avg/n497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18509.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18510 (.I0(\y_avg_black[6] ), .I1(n11675), .I2(n10838), 
            .O(\u_black_pixel_avg/n496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18510.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18511 (.I0(\y_avg_black[7] ), .I1(n11596), .I2(n10838), 
            .O(\u_black_pixel_avg/n495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18511.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18512 (.I0(\y_avg_black[8] ), .I1(n11538), .I2(n10838), 
            .O(\u_black_pixel_avg/n494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18512.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18513 (.I0(\y_avg_black[9] ), .I1(n11489), .I2(n10838), 
            .O(\u_black_pixel_avg/n493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18513.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18514 (.I0(\y_avg_black[10] ), .I1(n11448), .I2(n10838), 
            .O(\u_black_pixel_avg/n492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18514.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18515 (.I0(\y_avg_black[11] ), .I1(n11414), .I2(n10838), 
            .O(\u_black_pixel_avg/n491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18515.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18516 (.I0(\u_black_pixel_avg/x_sum[2] ), .I1(n4072), 
            .I2(n9701), .O(\u_black_pixel_avg/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18516.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18517 (.I0(\u_black_pixel_avg/x_sum[3] ), .I1(n4070), 
            .I2(n9701), .O(\u_black_pixel_avg/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18517.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18518 (.I0(\u_black_pixel_avg/x_sum[4] ), .I1(n4068), 
            .I2(n9701), .O(\u_black_pixel_avg/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18518.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18519 (.I0(\u_black_pixel_avg/x_sum[5] ), .I1(n4066), 
            .I2(n9701), .O(\u_black_pixel_avg/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18519.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18520 (.I0(\u_black_pixel_avg/x_sum[6] ), .I1(n4064), 
            .I2(n9701), .O(\u_black_pixel_avg/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18520.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18521 (.I0(\u_black_pixel_avg/x_sum[7] ), .I1(n4062), 
            .I2(n9701), .O(\u_black_pixel_avg/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18521.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18522 (.I0(\u_black_pixel_avg/x_sum[8] ), .I1(n4060), 
            .I2(n9701), .O(\u_black_pixel_avg/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18522.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18523 (.I0(\u_black_pixel_avg/x_sum[9] ), .I1(n4058), 
            .I2(n9701), .O(\u_black_pixel_avg/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18523.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18524 (.I0(\u_black_pixel_avg/x_sum[10] ), .I1(n4056), 
            .I2(n9701), .O(\u_black_pixel_avg/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18524.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18525 (.I0(\u_black_pixel_avg/x_sum[11] ), .I1(n4054), 
            .I2(n9701), .O(\u_black_pixel_avg/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18525.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18526 (.I0(\u_black_pixel_avg/x_sum[12] ), .I1(n4052), 
            .I2(n9701), .O(\u_black_pixel_avg/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18526.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18527 (.I0(\u_black_pixel_avg/x_sum[13] ), .I1(n4050), 
            .I2(n9701), .O(\u_black_pixel_avg/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18527.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18528 (.I0(\u_black_pixel_avg/x_sum[14] ), .I1(n4048), 
            .I2(n9701), .O(\u_black_pixel_avg/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18528.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18529 (.I0(\u_black_pixel_avg/x_sum[15] ), .I1(n4046), 
            .I2(n9701), .O(\u_black_pixel_avg/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18529.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18530 (.I0(\u_black_pixel_avg/x_sum[16] ), .I1(n4044), 
            .I2(n9701), .O(\u_black_pixel_avg/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18530.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18531 (.I0(\u_black_pixel_avg/x_sum[17] ), .I1(n4042), 
            .I2(n9701), .O(\u_black_pixel_avg/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18531.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18532 (.I0(\u_black_pixel_avg/x_sum[18] ), .I1(n4040), 
            .I2(n9701), .O(\u_black_pixel_avg/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18532.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18533 (.I0(\u_black_pixel_avg/x_sum[19] ), .I1(n4038), 
            .I2(n9701), .O(\u_black_pixel_avg/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18533.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18534 (.I0(\u_black_pixel_avg/x_sum[20] ), .I1(n4036), 
            .I2(n9701), .O(\u_black_pixel_avg/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18534.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18535 (.I0(\u_black_pixel_avg/x_sum[21] ), .I1(n4034), 
            .I2(n9701), .O(\u_black_pixel_avg/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18535.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18536 (.I0(\u_black_pixel_avg/x_sum[22] ), .I1(n4032), 
            .I2(n9701), .O(\u_black_pixel_avg/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18536.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18537 (.I0(\u_black_pixel_avg/x_sum[23] ), .I1(n4030), 
            .I2(n9701), .O(\u_black_pixel_avg/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18537.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18538 (.I0(\u_black_pixel_avg/x_sum[24] ), .I1(n4028), 
            .I2(n9701), .O(\u_black_pixel_avg/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18538.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18539 (.I0(\u_black_pixel_avg/x_sum[25] ), .I1(n4026), 
            .I2(n9701), .O(\u_black_pixel_avg/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18539.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18540 (.I0(\u_black_pixel_avg/x_sum[26] ), .I1(n4024), 
            .I2(n9701), .O(\u_black_pixel_avg/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18540.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18541 (.I0(\u_black_pixel_avg/x_sum[27] ), .I1(n4022), 
            .I2(n9701), .O(\u_black_pixel_avg/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18541.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18542 (.I0(\u_black_pixel_avg/x_sum[28] ), .I1(n4020), 
            .I2(n9701), .O(\u_black_pixel_avg/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18542.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18543 (.I0(\u_black_pixel_avg/x_sum[29] ), .I1(n4018), 
            .I2(n9701), .O(\u_black_pixel_avg/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18543.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18544 (.I0(\u_black_pixel_avg/x_sum[30] ), .I1(n4016), 
            .I2(n9701), .O(\u_black_pixel_avg/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18544.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18545 (.I0(\u_black_pixel_avg/x_sum[31] ), .I1(n4015), 
            .I2(n9701), .O(\u_black_pixel_avg/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18545.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18546 (.I0(\u_state_machine/current_state.WAITING ), .I1(\u_state_machine/current_state.WORKING ), 
            .O(\u_state_machine/equal_19/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__18546.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__18547 (.I0(\y_avg_black[4] ), .I1(\y_avg_black[3] ), .I2(\y_avg_black[5] ), 
            .I3(\y_avg_black[6] ), .O(n12102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__18547.LUTMASK = 16'he000;
    EFX_LUT4 LUT__18548 (.I0(\y_avg_black[9] ), .I1(\y_avg_black[10] ), 
            .I2(\y_avg_black[11] ), .O(n12103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__18548.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__18549 (.I0(\y_avg_black[7] ), .I1(n12102), .I2(\y_avg_black[8] ), 
            .I3(n12103), .O(n12104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__18549.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__18550 (.I0(\u_state_machine/equal_19/n3 ), .I1(n12104), 
            .I2(\u_state_machine/key0_debounced ), .O(n12105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__18550.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__18551 (.I0(\x_avg_black[6] ), .I1(\x_avg_black[7] ), .I2(\x_avg_black[9] ), 
            .I3(\x_avg_black[8] ), .O(n12106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h71cf */ ;
    defparam LUT__18551.LUTMASK = 16'h71cf;
    EFX_LUT4 LUT__18552 (.I0(\x_avg_black[10] ), .I1(\x_avg_black[11] ), 
            .I2(n12106), .O(n12107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__18552.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__18553 (.I0(\x_avg_black[8] ), .I1(\x_avg_black[7] ), .I2(\x_avg_black[9] ), 
            .O(n12108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__18553.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__18554 (.I0(n12108), .I1(\x_avg_black[10] ), .I2(\x_avg_black[11] ), 
            .O(n12109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__18554.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__18555 (.I0(n12107), .I1(n12109), .O(n12110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18555.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18556 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[0]), 
            .I2(n12105), .I3(n12110), .O(\u_state_machine/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__18556.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__18557 (.I0(\u_state_machine/counter_10s[4] ), .I1(\u_state_machine/counter_10s[5] ), 
            .I2(\u_state_machine/counter_10s[6] ), .I3(\u_state_machine/counter_10s[7] ), 
            .O(n12111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__18557.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__18558 (.I0(\u_state_machine/counter_10s[8] ), .I1(\u_state_machine/counter_10s[9] ), 
            .I2(\u_state_machine/counter_10s[10] ), .O(n12112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18558.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18559 (.I0(n12112), .I1(n12111), .I2(\u_state_machine/counter_10s[11] ), 
            .O(n12113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__18559.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__18560 (.I0(\u_state_machine/counter_10s[12] ), .I1(\u_state_machine/counter_10s[13] ), 
            .I2(\u_state_machine/counter_10s[14] ), .I3(\u_state_machine/counter_10s[15] ), 
            .O(n12114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__18560.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__18561 (.I0(n12114), .I1(n12113), .I2(\u_state_machine/counter_10s[16] ), 
            .I3(\u_state_machine/counter_10s[17] ), .O(n12115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__18561.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__18562 (.I0(n12115), .I1(\u_state_machine/counter_10s[18] ), 
            .I2(\u_state_machine/counter_10s[19] ), .O(n12116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__18562.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__18563 (.I0(\u_state_machine/counter_10s[20] ), .I1(n12116), 
            .I2(\u_state_machine/counter_10s[21] ), .I3(\u_state_machine/counter_10s[22] ), 
            .O(n12117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__18563.LUTMASK = 16'he000;
    EFX_LUT4 LUT__18564 (.I0(\u_state_machine/counter_10s[23] ), .I1(\u_state_machine/counter_10s[24] ), 
            .I2(\u_state_machine/counter_10s[25] ), .O(n12118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__18564.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__18566 (.I0(n12117), .I1(n12118), .I2(\u_state_machine/counter_10s[26] ), 
            .O(n12120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__18566.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__18567 (.I0(n12120), .I1(\u_state_machine/counter_10s[0] ), 
            .O(\u_state_machine/n99 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18567.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18568 (.I0(n12107), .I1(\u_state_machine/key0_debounced ), 
            .I2(zone_bit0), .I3(\u_state_machine/equal_19/n3 ), .O(\u_state_machine/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__18568.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__18569 (.I0(n12109), .I1(\u_state_machine/key0_debounced ), 
            .I2(zone_bit1), .I3(\u_state_machine/equal_19/n3 ), .O(\u_state_machine/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__18569.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__18570 (.I0(n12104), .I1(\u_state_machine/equal_19/n3 ), 
            .I2(\u_state_machine/key0_debounced ), .O(n12121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__18570.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__18571 (.I0(\u_state_machine/equal_19/n3 ), .I1(zone_bit2), 
            .I2(n12121), .O(\u_state_machine/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__18571.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__18572 (.I0(\u_state_machine/key0_debounced ), .I1(n12120), 
            .I2(\u_state_machine/equal_19/n3 ), .O(\u_state_machine/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__18572.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__18573 (.I0(\u_state_machine/key0_last ), .I1(key0), .O(\u_state_machine/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18573.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18574 (.I0(n12107), .I1(n12109), .O(n12122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18574.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18575 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[1]), 
            .I2(n12105), .I3(n12122), .O(\u_state_machine/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__18575.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__18576 (.I0(n12109), .I1(n12105), .O(n12123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18576.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18577 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[2]), 
            .I2(n12123), .I3(n12107), .O(\u_state_machine/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__18577.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__18578 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[3]), 
            .I2(n12107), .I3(n12123), .O(\u_state_machine/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__18578.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__18579 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[4]), 
            .I2(n12110), .I3(n12121), .O(\u_state_machine/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__18579.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__18580 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[5]), 
            .I2(n12121), .I3(n12122), .O(\u_state_machine/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__18580.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__18581 (.I0(n12109), .I1(n12121), .O(n12124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__18581.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__18582 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[6]), 
            .I2(n12124), .I3(n12107), .O(\u_state_machine/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__18582.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__18583 (.I0(\u_state_machine/equal_19/n3 ), .I1(led_data[7]), 
            .I2(n12107), .I3(n12124), .O(\u_state_machine/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__18583.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__18584 (.I0(n12120), .I1(\u_state_machine/counter_10s[0] ), 
            .O(n12125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18584.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18585 (.I0(n12125), .I1(\u_state_machine/counter_10s[1] ), 
            .O(\u_state_machine/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18585.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18586 (.I0(n12125), .I1(\u_state_machine/counter_10s[1] ), 
            .O(n12126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18586.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18587 (.I0(n12126), .I1(\u_state_machine/counter_10s[2] ), 
            .O(\u_state_machine/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18587.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18588 (.I0(n12126), .I1(\u_state_machine/counter_10s[2] ), 
            .O(n12127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18588.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18589 (.I0(n12127), .I1(\u_state_machine/counter_10s[3] ), 
            .O(\u_state_machine/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18589.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18590 (.I0(n12127), .I1(\u_state_machine/counter_10s[3] ), 
            .O(n12128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18590.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18591 (.I0(n12128), .I1(\u_state_machine/counter_10s[4] ), 
            .O(\u_state_machine/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18591.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18592 (.I0(n12128), .I1(\u_state_machine/counter_10s[4] ), 
            .O(n12129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18592.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18593 (.I0(n12129), .I1(\u_state_machine/counter_10s[5] ), 
            .O(\u_state_machine/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18593.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18594 (.I0(n12129), .I1(\u_state_machine/counter_10s[5] ), 
            .O(n12130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18594.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18595 (.I0(n12130), .I1(\u_state_machine/counter_10s[6] ), 
            .O(\u_state_machine/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18595.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18596 (.I0(n12130), .I1(\u_state_machine/counter_10s[6] ), 
            .I2(\u_state_machine/counter_10s[7] ), .O(\u_state_machine/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18596.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18597 (.I0(n12130), .I1(\u_state_machine/counter_10s[6] ), 
            .I2(\u_state_machine/counter_10s[7] ), .O(n12131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18597.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18598 (.I0(n12131), .I1(\u_state_machine/counter_10s[8] ), 
            .O(\u_state_machine/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18598.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18599 (.I0(n12130), .I1(\u_state_machine/counter_10s[6] ), 
            .I2(\u_state_machine/counter_10s[7] ), .I3(\u_state_machine/counter_10s[8] ), 
            .O(n12132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__18599.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__18600 (.I0(n12132), .I1(\u_state_machine/counter_10s[9] ), 
            .O(\u_state_machine/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18600.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18601 (.I0(n12132), .I1(\u_state_machine/counter_10s[9] ), 
            .I2(\u_state_machine/counter_10s[10] ), .O(\u_state_machine/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18601.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18602 (.I0(n12131), .I1(n12112), .I2(\u_state_machine/counter_10s[11] ), 
            .O(\u_state_machine/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18602.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18603 (.I0(n12131), .I1(n12112), .I2(\u_state_machine/counter_10s[11] ), 
            .O(n12133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18603.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18604 (.I0(n12133), .I1(\u_state_machine/counter_10s[12] ), 
            .O(\u_state_machine/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18604.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18605 (.I0(n12133), .I1(\u_state_machine/counter_10s[12] ), 
            .I2(\u_state_machine/counter_10s[13] ), .O(\u_state_machine/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18605.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18606 (.I0(\u_state_machine/counter_10s[12] ), .I1(\u_state_machine/counter_10s[13] ), 
            .I2(n12133), .O(n12134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18606.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18607 (.I0(n12134), .I1(\u_state_machine/counter_10s[14] ), 
            .O(\u_state_machine/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18607.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18608 (.I0(n12134), .I1(\u_state_machine/counter_10s[14] ), 
            .I2(\u_state_machine/counter_10s[15] ), .O(\u_state_machine/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18608.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18609 (.I0(n12131), .I1(n12112), .I2(n12114), .I3(\u_state_machine/counter_10s[11] ), 
            .O(n12135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__18609.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__18610 (.I0(n12135), .I1(\u_state_machine/counter_10s[16] ), 
            .O(\u_state_machine/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18610.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18611 (.I0(n12135), .I1(\u_state_machine/counter_10s[16] ), 
            .I2(\u_state_machine/counter_10s[17] ), .O(\u_state_machine/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18611.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18612 (.I0(n12135), .I1(\u_state_machine/counter_10s[16] ), 
            .I2(\u_state_machine/counter_10s[17] ), .O(n12136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18612.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18613 (.I0(n12136), .I1(\u_state_machine/counter_10s[18] ), 
            .O(\u_state_machine/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18613.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18614 (.I0(n12136), .I1(\u_state_machine/counter_10s[18] ), 
            .I2(\u_state_machine/counter_10s[19] ), .O(\u_state_machine/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18614.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18615 (.I0(n12136), .I1(\u_state_machine/counter_10s[18] ), 
            .I2(\u_state_machine/counter_10s[19] ), .O(n12137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__18615.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__18616 (.I0(n12137), .I1(\u_state_machine/counter_10s[20] ), 
            .O(\u_state_machine/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18616.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18617 (.I0(n12137), .I1(\u_state_machine/counter_10s[20] ), 
            .O(n12138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__18617.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__18618 (.I0(n12138), .I1(\u_state_machine/counter_10s[21] ), 
            .O(\u_state_machine/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18618.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18619 (.I0(n12138), .I1(\u_state_machine/counter_10s[21] ), 
            .I2(\u_state_machine/counter_10s[22] ), .O(\u_state_machine/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18619.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18620 (.I0(n12138), .I1(\u_state_machine/counter_10s[21] ), 
            .I2(\u_state_machine/counter_10s[22] ), .I3(\u_state_machine/counter_10s[23] ), 
            .O(\u_state_machine/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__18620.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__18621 (.I0(n12138), .I1(\u_state_machine/counter_10s[21] ), 
            .I2(\u_state_machine/counter_10s[22] ), .I3(\u_state_machine/counter_10s[23] ), 
            .O(n12139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__18621.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__18622 (.I0(n12139), .I1(\u_state_machine/counter_10s[24] ), 
            .O(\u_state_machine/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__18622.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__18623 (.I0(n12139), .I1(\u_state_machine/counter_10s[24] ), 
            .I2(\u_state_machine/counter_10s[25] ), .O(\u_state_machine/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__18623.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__18624 (.I0(n12139), .I1(\u_state_machine/counter_10s[24] ), 
            .I2(\u_state_machine/counter_10s[25] ), .I3(\u_state_machine/counter_10s[26] ), 
            .O(\u_state_machine/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80 */ ;
    defparam LUT__18624.LUTMASK = 16'hff80;
    EFX_LUT4 LUT__18625 (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(lcd_hs), .I2(\u_lcd_driver/r_lcd_dv ), 
            .O(\u_rgb2dvi/enc_0/n869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__18625.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__18626 (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(lcd_hs), .I2(\u_lcd_driver/r_lcd_dv ), 
            .O(\u_rgb2dvi/enc_0/n770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__18626.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__18627 (.I0(\u_lcd_driver/r_lcd_rgb[23] ), .I1(lcd_hs), 
            .I2(\u_lcd_driver/r_lcd_dv ), .O(\u_rgb2dvi/enc_0/n806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__18627.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__18628 (.I0(lcd_hs), .I1(lcd_vs), .O(n12140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__18628.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__18629 (.I0(n12140), .I1(\u_lcd_driver/r_lcd_rgb[23] ), 
            .I2(\u_rgb2dvi/enc_0/acc[4] ), .I3(\u_lcd_driver/r_lcd_dv ), 
            .O(\u_rgb2dvi/enc_0/n812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__18629.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__18630 (.I0(\r_hdmi_tx0_o[6] ), .I1(\w_hdmi_txd0[0] ), 
            .I2(rc_hdmi_tx), .O(n926_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18630.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18631 (.I0(\r_hdmi_tx0_o[7] ), .I1(\w_hdmi_txd0[4] ), 
            .I2(rc_hdmi_tx), .O(n925_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18631.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18632 (.I0(\r_hdmi_tx0_o[8] ), .I1(\w_hdmi_txd0[0] ), 
            .I2(rc_hdmi_tx), .O(n924_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18632.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18633 (.I0(\r_hdmi_tx0_o[9] ), .I1(\w_hdmi_txd0[4] ), 
            .I2(rc_hdmi_tx), .O(n923_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18633.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18634 (.I0(\r_hdmi_tx1_o[6] ), .I1(\w_hdmi_txd1[0] ), 
            .I2(rc_hdmi_tx), .O(n937_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18634.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18635 (.I0(\r_hdmi_tx1_o[7] ), .I1(\w_hdmi_txd1[4] ), 
            .I2(rc_hdmi_tx), .O(n936_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18635.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18636 (.I0(\r_hdmi_tx1_o[8] ), .I1(\w_hdmi_txd1[0] ), 
            .I2(rc_hdmi_tx), .O(n935_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18636.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18637 (.I0(\r_hdmi_tx1_o[9] ), .I1(\w_hdmi_txd1[4] ), 
            .I2(rc_hdmi_tx), .O(n934_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18637.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18638 (.I0(\r_hdmi_tx2_o[6] ), .I1(\w_hdmi_txd2[0] ), 
            .I2(rc_hdmi_tx), .O(n948_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18638.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18639 (.I0(\r_hdmi_tx2_o[7] ), .I1(\w_hdmi_txd2[4] ), 
            .I2(rc_hdmi_tx), .O(n947_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18639.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18640 (.I0(\r_hdmi_tx1_o[8] ), .I1(\w_hdmi_txd2[0] ), 
            .I2(rc_hdmi_tx), .O(n946_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__18640.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__18641 (.I0(\r_hdmi_tx2_o[9] ), .I1(\w_hdmi_txd2[4] ), 
            .I2(rc_hdmi_tx), .O(n945_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__18641.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__18642 (.I0(n1735), .I1(\PowerOnResetCnt[1] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n32_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__18642.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__18643 (.I0(n1733), .I1(\PowerOnResetCnt[2] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n31_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__18643.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__18644 (.I0(n1731), .I1(\PowerOnResetCnt[3] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n30_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__18644.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__18645 (.I0(n1729), .I1(\PowerOnResetCnt[4] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n29_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__18645.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__18646 (.I0(n1727), .I1(\PowerOnResetCnt[5] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n28_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__18646.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__18647 (.I0(n1725), .I1(\PowerOnResetCnt[6] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n27_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__18647.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__18648 (.I0(n1724), .I1(\PowerOnResetCnt[7] ), .I2(hdmi_resetn_o), 
            .I3(PllLocked[0]), .O(n26_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__18648.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__18784 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
            .O(DdrCtrl_CFG_SEQ_RST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__18784.LUTMASK = 16'h5555;
    EFX_GBUFCE CLKBUF__3 (.CE(1'b1), .I(hdmi_clk1x_i), .O(\hdmi_clk1x_i~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__3.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__2 (.CE(1'b1), .I(Axi0Clk), .O(\Axi0Clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__2.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(cmos_pclk), .O(\cmos_pclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(hdmi_clk2x_i), .O(\hdmi_clk2x_i~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2  (.I0(n3493), .I1(1'b1), 
            .CI(1'b0), .CO(n12216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(79)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2  (.I0(n3493), .I1(1'b1), 
            .CI(1'b0), .CO(n12215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(1'b0), .I1(1'b0), 
            .CI(n12214), .O(n3493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n12213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n12212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\hdmi_ip\tmds_channel.v(93)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2952/i5  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2952/i5 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2952/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2876/i6  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2876/i6 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2876/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2798/i7  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2798/i7 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2798/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2718/i8  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2718/i8 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2718/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2636/i9  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2636/i9 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2636/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2552/i10  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2552/i10 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2552/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2466/i11  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2466/i11 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2466/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2378/i12  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2378/i12 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2378/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2288/i13  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2288/i13 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2288/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2196/i14  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2196/i14 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2196/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2102/i15  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2102/i15 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2102/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2006/i16  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2006/i16 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_2006/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1908/i17  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1908/i17 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1908/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1808/i18  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1808/i18 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1808/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1706/i19  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1706/i19 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1706/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1602/i20  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1602/i20 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1602/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1496/i21  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1496/i21 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1496/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1388/i22  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1388/i22 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1388/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1278/i23  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1278/i23 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1278/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1166/i24  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1166/i24 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1166/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1052/i25  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1052/i25 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_1052/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_936/i26  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_936/i26 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_936/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_818/i27  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_818/i27 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_818/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_698/i28  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_698/i28 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_698/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_576/i29  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_576/i29 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_576/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_452/i30  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_452/i30 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_452/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_326/i31  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_326/i31 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_326/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_24/add_198/i32  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(48)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_198/i32 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_24/add_198/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2718/i8  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2718/i8 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2718/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2636/i9  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2636/i9 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2636/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2552/i10  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2552/i10 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2552/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2466/i11  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2466/i11 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2466/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2378/i12  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2378/i12 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2378/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2288/i13  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2288/i13 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2288/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2196/i14  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2196/i14 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2196/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2102/i15  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2102/i15 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2102/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2006/i16  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2006/i16 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_2006/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1908/i17  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1908/i17 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1908/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1808/i18  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1808/i18 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1808/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1706/i19  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1706/i19 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1706/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1602/i20  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1602/i20 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1602/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1496/i21  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1496/i21 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1496/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1388/i22  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1388/i22 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1388/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1278/i23  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1278/i23 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1278/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1166/i24  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1166/i24 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1166/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1052/i25  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1052/i25 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_1052/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_936/i26  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_936/i26 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_936/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_818/i27  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_818/i27 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_818/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_698/i28  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_698/i28 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_698/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_576/i29  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_576/i29 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_576/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_452/i30  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_452/i30 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_452/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_326/i31  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_326/i31 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_326/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_black_pixel_avg/div_23/add_198/i32  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\black_pixel_avg.v(47)
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_198/i32 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_black_pixel_avg/div_23/add_198/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_lcd_driver/sub_61/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n12149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(148)
    defparam \AUX_ADD_CI__u_lcd_driver/sub_61/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_lcd_driver/sub_61/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(167)
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl_0/sub_131/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n12144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\axi\axi4_ctrl.v(356)
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/sub_131/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/sub_131/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_R0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1279)
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_56/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n12142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Efinity\ip\W0_FIFO_128\W0_FIFO_128.v(1277)
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl_0/u_W0_FIFO_128/u_efx_fifo_top/xefx_fifo_ctl/sub_53/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_lcd_driver/sub_60/add_2/i2  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n12148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\code\learning\a241111_03\Source\lcd_driver.v(147)
    defparam \AUX_ADD_CI__u_lcd_driver/sub_60/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_lcd_driver/sub_60/add_2/i2 .I1_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_14282319_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_14282319_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_14282319_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_14282319_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_14282319_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__16_16_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__16_16_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__16_16_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__16_16_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__16_16_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__20_20_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_14282319__16_16_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_14282319_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_237
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_238
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_239
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_240
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_241
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_242
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_243
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_244
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_245
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_246
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_247
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_248
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_249
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_250
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_251
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_252
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_253
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_254
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_255
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_256
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_257
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_258
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_259
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_260
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_261
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_262
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_263
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_264
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_265
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_266
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_267
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_268
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_269
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_270
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_271
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_272
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_273
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_274
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_275
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_276
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_277
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_278
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_279
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_14282319_280
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_14282319_0
// module not written out since it is a black box. 
//

